library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;
use IEEE.NUMERIC_STD.ALL;
entity coefficient_memory is
  generic(
    data : integer := 16;
    addr_data : integer := 15
    );
  port ( 
    CLK : in std_logic;
    ADDRESS_DATA,RESET_ADDRESS : in std_logic_vector(addr_data-1 downto 0); --address of operand
    DATA_RAM_IN,RESET_DATA : in std_logic_vector(data-1 downto 0); --value of operand
    DATA_RAM_OUT : out std_logic_vector(data-1 downto 0);
    READ_RAM,WRITE_RAM,WRITE_RESET : in std_logic --read and write operation 
    );
end coefficient_memory;

architecture Behavioral of coefficient_memory is
type ram is array (0 to 32767) of integer;
signal RAM_DATA : ram := ( 
-- gaussian approx - 20x16
/*

--RVFL 16


-78,52,64,85,75,70,68,457,66,64,38,4461,0,67,-1,101,10,133,6,250,
0,58,27,56,-50,67,-74,61,-76,358,9,1022,-67,4899,74,1824,75,94,-19,72,
-1,55,8,86,-41,69,24,53,-20,110,-32,77,47,16711,3,229,-31,70,-51,60,
-59,1955,32,280,60,349,22,273,-48,408,75,173,41,54,64,53,-26,84,62,158,
-57,319,-18,84,65,75,-6,160,-25,61,-44,59,-38,154,-40,75,37,78,-67,125,
-45,104,31,928,41,54,-72,74,-9,59,-58,150,-64,168,3,51,32,82,49,50,
-13,68,52,67,-24,1542,-74,632,0,435,18,54,67,184,1,135,36,133,29,197,
-40,140,-5,248,-6,270,-53,1527,-14,69,-1,380,3,203,50,65,63,153,-6,66,
-67,88,70,55,18,65,47,153,-46,54,-51,91,-59,64,-68,83,35,89,26,123,
-25,1099,49,105,-1,1194,-54,129,-45,129,-63,169,-62,189,54,83,29,66,-35,158,
-53,78,77,113,-4,179,-58,91,-43,64,6,62,55,69,49,441,55,54,58,64,
61,73,-53,367,-10,58,-24,90,37,54,-34,148,7,74,-15,225,23,60,-51,111,
72,126,3,61,59,135,-2,151,-13,10098,-64,413,-38,90,-74,691,-32,90,13,70,
-74,365,71,54,-50,55,32,117,13,183,-2,109,12,73,43,98,53,60,-6,225,
32,120,24,71,30,172,48,198,-1,1369,21,200,-30,287,29,144,-41,1771,28,60,
12,67,58,74,33,131,-37,246,-11,251,-74,67,47,107,67,254,33,62,-4,69,


-181,-73,21,-95,573,-50,291,93,137,-331,-13,-177,94,70,-363,-39,
32,140,-52,-423,22,-666,-510,162,819,-127,474,-596,285,18,-294,360,
-335,-172,-348,-109,-38,-54,113,-628,217,249,58,397,716,390,-247,-240,
104,63,-172,422,66,-145,-62,89,-267,166,-188,115,80,-191,280,-44,
498,13,642,236,-1279,-1,187,-390,-938,935,-154,671,-118,364,-32,-361,
72,-88,19,-431,-135,161,205,-194,248,-96,-7,-168,-38,346,74,-135,
1,-102,387,289,418,-178,-232,240,92,215,-71,309,-774,-660,132,136,
-302,-128,35,203,-53,-462,-377,-334,767,903,4,298,120,-558,-169,252,
46,17,-442,81,349,-411,-146,-184,686,542,-127,95,-277,-253,-151,202,
276,53,-129,-26,-234,443,480,370,-640,-872,-147,-246,71,455,227,-173,
-102,9,-210,51,-166,1135,74,241,-615,-462,-35,529,-201,-598,525,-14,
-126,-33,-206,-37,300,429,313,-183,-1167,-385,334,-87,545,645,194,-473,
-29,274,259,-108,564,19,-216,305,-377,-289,22,-300,-474,-181,35,492,
-129,129,74,123,-501,125,-140,-21,615,-482,97,-232,-223,247,-138,4,
16,-68,-74,-211,-110,132,56,188,397,260,-79,-614,322,127,-178,-56,

*/
/*
--RVFL 32
-78,100,75,58,66,82,0,101,10,84,72,66,33,1394,44,103,38,322,-20,120,
0,63,-50,138,-76,74,-67,93,75,363,57,2968,39,128,-58,158,-78,75,4,914,
-1,54,-41,60,-20,245,47,53,-31,84,64,116,34,52,-8,294,-80,64,34,8202,
-59,63,60,191,-48,155,41,129,-26,60,-76,62,-57,350,-60,715,67,5388,14,64,
-57,167,65,50,-25,51,-38,95,37,122,-55,337,27,135,51,246,-28,78,22,56,
-45,69,41,125,-9,182,-64,258,32,870,-4,66,66,53,55,122,-33,93,17,169,
-13,81,-24,90,0,71,67,1485,36,223,38,143,-75,5947,-62,75,-37,381,-20,124,
-40,59,-6,77,-14,188,3,96,63,88,-23,1160,-50,59,35,188,-41,589,-28,53,
-67,123,18,159,-46,87,-59,500,35,81,10,69,42,59,68,56,44,52,10,125,
-25,110,-1,57,-45,57,-62,73,29,52,-73,58,-73,63,-18,722,-38,52,40,101,
-53,533,-4,50,-43,61,55,214,55,55,22,51,-35,56,44,62,35,156,67,741,
61,228,-10,87,37,1710,7,98,23,171,29,328,57,131,68,106,28,126,52,98,
72,94,59,224,-13,117,-38,61,-32,437,-17,84,-21,168,-79,157,8,450,9,70,
-74,94,-50,174,13,127,12,72,53,60,-58,183,64,95,-36,355,29,200,52,178,
32,70,30,61,-1,55,-30,117,-41,95,-13,56,-34,170,-74,83,-52,154,-75,108,
12,174,33,89,-11,1396,47,73,33,51,38,546,-19,202,-48,87,-6,72,48,822,
64,430,68,92,38,109,-1,155,6,716,13,276,-63,810,-78,72,-1,116,-48,82,
27,267,-74,334,9,50,74,54,-19,142,61,638,50,141,-72,58,-76,80,30,70,
8,115,24,67,-32,1373,3,161,-51,67,13,168,69,318,24,108,-45,76,52,2127,
32,269,22,319,75,74,64,81,62,88,-52,52,-51,65,-34,52,69,94,-30,104,
-18,404,-6,267,-44,68,-40,112,-67,61,15,136,-30,73,55,50,25,92,-16,582,
31,68,-72,85,-58,476,3,961,49,67,-71,89,28,57,-27,420,77,32767,78,51,
52,54,-74,80,18,191,1,123,29,140,39,126,-67,104,67,91,-21,78,-39,115,
-5,820,-53,263,-1,105,50,84,-6,130,-48,50,-75,205,-59,83,42,72,41,100,
70,1195,47,53,-51,248,-68,105,26,219,65,69,-28,65,8,3348,16,50,-15,101,
49,175,-54,70,-63,53,54,53,-35,61,-4,59,-18,262,-33,339,16,107,-30,53,
77,86,-58,62,6,69,49,390,58,114,-9,392,8,130,49,67,-62,73,43,78,
-53,53,-24,64,-34,494,-15,66,-51,59,-58,53,8,80,-26,134,-44,118,-8,68,
3,85,-2,95,-64,57,-74,80,13,52,49,182,-27,78,-61,61,-68,235,34,84,
71,73,32,79,-2,173,43,140,-6,146,67,72,-12,103,-7,50,1,353,-44,95,
24,76,48,2668,21,123,29,90,28,136,31,168,-40,78,-40,85,-25,552,52,61,
58,52,-37,85,-74,80,67,385,-4,104,27,77,-48,237,39,2407,-49,224,35,59,


-9,140,21,152,-75,414,-11,-350,-217,-3,-111,-367,-593,293,-68,84,-78,-148,-59,-89,-236,-124,-88,63,140,153,407,303,43,181,510,-332,
3,-139,340,-168,1106,-954,-137,-518,609,-562,148,264,371,262,673,-15,221,-151,-4,-125,27,-90,-46,-607,-596,-126,-782,-4,796,465,-489,84,
-87,-1,-329,-6,-679,178,-33,-241,189,576,-7,-3,-270,-379,-492,-44,-187,128,588,8,52,-93,-567,-674,-159,646,441,779,-922,325,922,22,
-38,-73,374,60,-204,-300,119,248,480,322,-239,-177,372,247,123,-154,639,168,197,-278,152,122,404,138,-407,-482,-263,-77,-451,168,-442,-138,
162,33,985,141,109,85,2,-168,-704,396,-135,634,450,-107,-543,413,-86,-52,-255,453,-113,165,-304,50,117,-1145,190,-631,-331,580,-614,109,
-277,114,-624,10,1,518,386,10,8,475,36,-135,-587,-163,-384,247,-498,314,-185,-234,25,-178,20,129,-305,424,326,-286,45,427,-19,161,
251,-98,481,86,343,-493,-244,-417,-485,-348,26,-204,131,264,115,-171,-87,-213,-58,107,227,233,1086,621,43,-946,-128,376,281,-185,-252,-187,
39,50,-271,-97,-166,238,188,204,371,255,109,148,167,-287,-722,-69,-49,-116,-213,-27,-488,22,44,-132,-134,559,129,-13,-424,-159,464,39,
-396,-18,-28,-52,54,-222,90,54,644,-75,13,-144,-343,-13,149,140,233,44,15,364,-198,-237,442,-188,-287,-119,-182,254,-427,361,54,-152,
48,108,-271,-86,62,275,-175,-39,-648,-327,124,195,-60,-266,-180,-136,42,-217,-15,761,-475,12,-162,-186,889,125,40,-14,440,-589,298,173,
-372,-142,-440,-82,110,-191,-123,-251,316,-47,64,-87,-253,294,1297,-246,92,214,-71,15,-357,96,308,79,-72,-241,171,344,179,-420,-287,119,
535,141,452,147,170,-9,24,-526,-94,400,60,153,210,-507,-349,-80,270,-306,70,-127,-249,119,-555,84,21,-562,100,-446,680,56,-2,-40,
275,-73,-54,19,-524,440,117,1602,-291,93,-95,-83,306,11,1135,-17,-327,154,-96,-557,708,-26,-237,114,399,675,-343,-1156,-82,-898,-70,-363,
-571,-76,-244,-29,-257,-163,-127,289,264,-261,-2,-291,-191,-24,-321,-25,273,158,105,39,182,-145,-207,671,128,262,-192,815,176,-172,-39,227,
484,20,-294,-77,-40,157,-102,170,-152,-415,30,24,294,32,-571,151,-401,100,20,-400,673,139,-194,-1,219,691,174,-345,-322,-192,-12,247,
*/

/*
--RVFL 64

-78,84,66,194,10,351,33,53,38,72,0,260,18,3332,15,76,-74,194,-55,62,
0,96,-76,160,75,59,39,90,-78,80,47,234,27,56,-58,60,-18,165,26,506,
-1,121,-20,219,-31,116,34,216,-80,82,67,199,-47,120,14,61,72,70,43,1758,
-59,97,-48,755,-26,91,-57,334,67,65,46,500,-29,212,53,205,-57,53,-79,80,
-57,866,-25,70,37,73,27,62,-28,188,-32,386,76,353,-15,261,-21,624,22,180,
-45,186,-9,95,32,86,66,561,-33,60,35,67,-36,50,-71,163,69,73,6,82,
-13,62,0,205,36,60,-75,203,-37,166,18,86,32,123,-44,107,-79,92,-59,60,
-40,53,-14,511,63,74,-50,54,-41,55,55,57,-38,81,11,324,54,288,-66,70,
-67,4165,-46,133,35,52,42,339,44,152,-15,2052,12,271,18,277,54,62,73,138,
-25,2953,-45,75,29,196,-73,81,-38,200,-7,92,60,1126,72,137,45,77,73,78,
-53,53,-43,146,55,79,-35,102,35,64,-65,62,51,159,64,56,61,101,-29,60,
61,59,37,120,23,81,57,463,28,441,-45,82,-75,136,-33,524,-19,87,-17,95,
72,101,-13,106,-32,71,-21,71,8,65,5,217,-12,69,-62,73,-32,384,-62,187,
-74,53,13,114,53,223,64,60,29,95,5,3011,-17,4000,51,78,4,61,-40,52,
32,199,-1,119,-41,664,-34,56,-52,76,34,68,64,53,4,63,-33,73,-28,268,
12,158,-11,132,33,2355,-19,219,-6,117,-34,62,-74,80,74,4117,-41,54,31,248,
64,53,38,137,6,107,-63,127,-1,128,-61,794,-7,399,-69,133,-70,144,-11,152,
27,148,9,71,-19,86,50,573,-76,54,-50,110,77,55,-24,64,-23,86,20,1450,
8,51,-32,66,-51,1475,69,55,-45,77,-11,166,-74,490,39,84,-55,563,25,73,
32,353,75,147,62,93,-51,500,69,184,-50,104,27,68,10,115,42,273,5,265,
-18,82,-44,64,-67,86,-30,55,25,334,-60,65,38,60,51,54,29,199,6,60,
31,82,-58,100,49,711,28,893,77,1691,36,88,-63,72,39,854,58,175,-80,377,
52,310,18,110,29,56,-67,127,-21,79,66,130,-38,250,-23,293,-3,150,22,53,
-5,246,-1,54,-6,467,-75,130,42,124,-70,71,-4,148,-19,488,-41,149,31,75,
70,122,-51,90,26,249,-28,96,16,71,-73,84,-48,515,-44,69,42,273,78,119,
49,99,-63,76,-35,139,-18,106,16,183,-34,57,69,95,49,70,-50,155,-6,384,
77,150,6,219,58,79,8,61,-62,62,13,286,35,106,-10,57,-19,54,29,93,
-53,74,-34,144,-51,146,8,65,-44,54,70,110,-64,66,55,56,20,78,-13,112,
3,52,-64,105,13,91,-27,72,-68,72,13,80,60,116,72,67,22,69,-46,58,
71,58,-2,81,-6,90,-12,55,1,110,29,147,-34,83,-25,387,-3,83,-57,111,
24,286,21,68,28,169,-40,1247,-25,90,24,85,-15,220,-21,99,22,228,-66,802,
58,98,-74,59,-4,136,-48,85,-49,274,71,713,19,241,-3,114,-46,54,-44,70,
75,50,0,71,72,55,44,111,-20,294,57,502,-1,460,40,266,-3,57,-14,83,
-50,107,-67,81,57,143,-58,51,4,784,-22,105,6,297,-77,96,-30,76,-71,92,
-41,57,47,103,64,55,-8,404,34,72,52,92,71,2102,-11,67,-53,50,-79,248,
60,619,41,120,-76,51,-60,228,14,177,-38,50,-18,130,48,106,-69,83,44,100,
65,71,-38,63,-55,64,51,105,22,51,78,75,3,50,-56,53,-48,1590,62,61,
41,317,-64,103,-4,109,55,613,17,66,-16,72,-49,59,41,55,-15,127,-33,80,
-24,54,67,288,38,52,-62,142,-20,73,9,80,-75,53,-24,79,26,70,-16,67,
-6,124,3,197,-23,228,35,164,-28,74,24,50,3,118,-73,112,-38,78,68,73,
18,121,-59,206,10,54,68,64,10,82,-30,58,-64,54,36,261,61,177,-16,177,
-1,524,-62,61,-73,63,-18,92,40,438,59,51,28,80,57,69,-69,232,-2,69,
-4,654,55,50,22,81,44,1535,67,51,78,62,-43,344,76,64,49,189,-69,50,
-10,81,7,62,29,58,68,75,52,94,11,86,1,129,-56,99,-5,54,1,99,
59,92,-38,69,-17,144,-79,64,9,74,-44,63,50,144,15,67,-29,105,34,146,
-50,143,12,83,-58,360,-36,53,52,82,-34,85,31,496,-36,61,-58,60,-35,5005,
30,51,-30,130,-13,4583,-74,61,-75,96,51,127,-12,394,61,66,15,221,-6,3004,
33,113,47,70,38,132,-48,72,48,184,10,208,29,75,-65,57,11,104,-70,493,
68,72,-1,92,13,115,-78,268,-48,82,7,82,-29,96,-51,97,30,127,17,132,
-74,210,74,148,61,68,-72,54,30,70,-56,458,66,239,-67,130,57,80,33,86,
24,99,3,607,13,293,24,350,52,134,38,65,-30,4366,-33,50,-6,138,-76,90,
22,53,64,240,-52,121,-34,56,-30,70,-55,139,18,111,72,54,72,51,-4,58,
-6,122,-40,51,15,106,55,97,-16,368,-50,50,-9,59,-21,55,78,105,-66,146,
-72,92,3,147,-71,57,-27,63,78,70,14,142,-72,51,10,58,-61,112,77,75,
-74,168,1,69,39,187,67,128,-39,64,19,59,-15,92,-17,510,7,174,-11,125,
-53,154,50,104,-48,95,-59,62,41,50,-50,69,14,57,77,122,16,57,0,143,
47,127,-68,85,65,612,8,86,-15,67,70,253,-4,58,34,233,-78,84,-1,304,
-54,195,54,176,-4,233,-33,121,-30,52,33,1220,70,201,55,1485,-56,1157,69,55,
-58,64,49,77,-9,239,49,129,43,206,48,150,-59,51,-60,96,39,72,23,89,
-24,98,-15,566,-58,133,-26,54,-8,59,45,63,40,89,70,68,-20,130,37,621,
-2,52,-74,77,49,66,-61,58,34,72,4,79,20,81,-36,160,50,111,15,52,
32,86,43,57,67,95,-7,94,-44,56,21,106,-23,51,30,115,79,118,3,62,
48,69,29,55,31,137,-40,184,52,638,-77,110,8,158,-32,167,14,123,51,91,
-37,107,67,83,27,124,39,92,35,90,13,89,-59,51,24,103,-77,57,54,90,

690,-477,-94,-179,29,-79,-310,979,216,7,-1416,-101,-368,-1056,-1577,-125,-287,-250,-159,43,871,-17,131,260,-437,235,46,254,587,990,-417,-201,416,-1355,70,318,426,955,798,-282,129,-539,386,-433,-319,184,-278,1374,233,-132,-744,21,-319,-221,826,-495,21,49,-727,475,-1479,1160,-225,600,
395,453,129,125,342,-296,631,389,-177,-279,1237,65,-307,207,894,-33,1577,-385,-1185,113,855,-124,-360,927,364,90,-874,94,2201,-1595,-338,2,91,353,-142,-944,-117,27,401,841,352,-127,-303,266,-1226,1477,-146,-387,143,-294,-43,541,-292,-176,-578,-870,-144,-152,-138,-310,-2009,224,-225,55,
-902,-102,-307,-553,-423,69,895,378,-424,-277,-121,15,594,1099,312,116,-416,90,1264,-91,-897,-41,-1025,865,201,191,-528,194,-2285,41,883,361,-393,1071,-156,-282,-553,34,290,485,-907,-330,-76,541,942,-1656,939,194,-1238,1064,-43,-1338,1336,-230,-1169,648,-326,418,659,839,1089,7,152,-266,
277,-497,218,713,347,-287,-290,618,-98,139,-474,393,-2140,-182,1045,35,732,-36,-287,-174,-431,221,245,118,136,494,550,-998,-29,20,39,-9,-107,342,-72,-983,376,356,1243,-442,-461,292,50,179,517,296,429,547,-1004,30,-1107,377,-501,90,230,-508,539,-37,-457,175,-215,158,-154,-165,
238,-525,-274,-65,51,126,74,-548,202,35,517,-301,627,246,93,-44,-325,-313,287,264,854,106,-35,-870,-396,1215,-354,-497,-418,517,-187,181,115,355,-26,72,47,336,-52,131,-3,-648,-14,-104,2,-27,-196,-934,-438,-127,10,-2,-279,26,691,339,-303,-93,519,44,407,-124,412,-650,
-196,609,430,300,-451,400,160,-824,-402,-124,-862,330,-914,-1269,-1057,-26,924,31,391,485,249,158,-49,-166,-76,-483,-148,259,822,-484,-943,-238,-108,16,-54,-137,524,-19,-292,514,745,447,-13,564,-20,264,568,886,44,1186,442,215,0,57,-47,155,0,59,-884,-647,-754,-606,-66,412,
257,-160,-254,249,156,-423,79,-689,755,105,1445,14,444,604,396,-13,-1534,-114,-525,118,49,-332,-303,-913,61,757,-490,52,331,1195,-368,242,-131,323,138,576,-343,-405,-475,-307,-229,-105,493,105,-259,-278,-754,-730,293,-1646,523,603,-1142,-172,1030,-466,111,-174,543,-150,1249,-60,-450,-65,
-325,-140,383,187,575,-657,-1757,-474,200,370,246,528,-528,-306,803,62,-18,1247,223,625,-1500,65,944,-239,500,-1446,1287,127,-259,-487,535,-506,-96,-602,110,-167,792,-1435,172,-620,-385,1410,-636,-25,432,705,-95,-762,1199,-1075,-647,-170,796,652,599,-251,284,-38,136,-101,1042,-643,334,-1090,
178,-149,160,530,188,252,301,-610,472,-33,-724,-312,-131,-110,-400,-8,538,-378,-358,-464,268,-89,264,339,89,253,-275,-845,-50,192,775,311,-101,-190,-46,-357,407,276,648,-650,472,-568,-2,132,1463,231,131,75,-950,705,139,-895,1711,-266,-526,646,-524,-122,43,-184,266,-733,-50,-472,
-241,356,-273,-698,-537,617,203,-700,234,-286,397,-707,2967,531,-586,-18,-874,-603,558,-32,616,-182,272,-569,-205,-255,-412,562,-473,240,-185,28,145,-529,40,1353,-1102,29,-1456,420,84,-596,236,-265,-340,-914,-494,-834,1136,302,1417,-650,1186,64,-302,813,-258,63,426,-240,430,-311,221,-40,
-201,78,83,115,69,-6,-145,-103,197,-51,808,-230,-318,200,445,22,440,-297,-98,-290,198,-9,-274,146,283,230,-244,-390,9,-112,-276,58,15,168,18,-108,-253,374,397,-49,-96,91,99,594,144,-287,-34,-7,0,-417,-42,-123,-214,163,-78,-260,-53,-98,-310,13,101,222,-139,-325,
-187,-689,55,-317,-122,274,291,-108,-46,-4,212,-244,-20,-861,-406,7,242,286,287,192,453,-10,-73,-555,-2,700,297,40,-1112,862,12,-146,20,-2,-78,242,-22,-85,-307,-286,-267,-90,190,235,-482,-3,252,-283,18,395,334,209,-332,794,436,-225,38,-54,-55,104,-1005,698,34,269,
-71,460,16,104,-206,331,312,682,-464,262,-1189,148,122,-217,-814,10,-101,736,-566,-1038,-478,27,431,391,-237,-742,815,-127,639,-109,780,121,-9,-401,66,588,494,-585,-825,-877,805,-389,34,-809,102,376,-32,314,-248,386,179,694,-541,-321,-649,587,129,62,117,-166,-105,-354,89,1079,
208,187,-55,-193,-30,109,145,925,-142,-26,-564,-363,-208,659,292,31,153,-197,117,-503,-635,125,142,815,-165,-429,235,-162,-428,-378,394,76,72,-14,9,-442,-168,607,-21,73,151,264,-378,-934,322,-287,199,49,-172,624,-479,-507,480,-46,-793,497,-61,16,419,141,210,111,122,214,
-215,558,-206,-284,-29,-419,-796,-119,-502,114,761,716,99,311,623,-14,-1036,143,188,687,-322,126,-298,-521,-174,-885,187,1281,384,-1022,-552,-253,98,498,127,161,-481,-369,-443,834,-432,969,122,177,-1208,-155,-487,501,955,-982,113,1177,-1709,-444,393,-679,566,91,-219,-39,734,126,-84,362,
*/






--MLP 16

-19,-141,-35,65,67,-59,20,47,-204,258,
-51,5,-23,-11,47,53,56,-47,0,-8,
18,35,-6,2,-101,-31,63,61,173,-196,
-3,-38,-97,-95,-45,135,-117,109,-121,122,
142,-21,4,-9,-9,-165,5,-9,-13,-5,
-153,49,34,-81,0,-53,2,-130,-28,53,
2,10,-12,18,1,-2,-22,14,16,10,
-46,111,88,139,-95,21,8,-29,-106,-14,
84,113,-41,-11,69,43,-20,-28,-124,-169,
-1,-20,0,-1,-20,-20,-21,-21,0,-1,
28,16,-107,-39,17,128,6,45,15,165,
52,-125,118,-121,24,126,-69,-60,-26,105,
-93,51,25,-174,148,-67,-101,9,99,-58,
6,6,6,1,24,4,14,-6,15,6,
-199,5,-85,113,20,-32,95,5,-32,-129,
327,-159,82,-72,-28,-42,56,-96,-14,-5,

-97,40,-220,2224,677,3487,125,-836,793,108,462,-659,2145,200,2802,-487,


-120,36,42,109,-106,-121,-40,29,45,-10,-23,-124,-136,-29,-116,115,-16,
-43,-40,-26,138,-95,187,-39,-24,-36,-11,-33,23,-67,-42,-105,127,-26,
34,-2,-75,162,-92,-165,-13,-27,-9,-10,-27,-94,123,-33,-67,-85,-3,
97,7,-85,159,-40,0,-78,-132,-41,-19,-10,-202,21,-68,114,128,-53,
-9,38,-16,-59,-109,-106,-8,-4,22,-20,-18,58,14,-28,-94,54,-8,
-64,-47,-12,-118,54,110,-56,-60,46,20,-34,-120,84,-37,31,55,-22,
-148,62,-13,17,117,-146,-66,3,-116,0,-21,41,60,-48,-121,102,-38,
-160,33,6,-98,-149,-80,-3,-19,-106,-10,10,-99,53,-3,108,28,5,
31,-143,-87,-28,-78,-25,-11,2,-83,0,92,-8,-43,-32,-5,45,-2,
-139,-77,83,68,13,73,-51,129,86,-1,-71,57,24,-53,98,-179,-42,
21,44,35,-45,-40,-37,-11,-2,32,20,-2,2,-59,-21,3,-62,-2,
56,-33,104,6,10,-9,-35,-7,-40,-10,-17,-10,-29,-37,-45,-10,-14,
111,87,-57,-39,-106,13,-28,-1,-66,0,-10,-138,-21,-28,-66,32,-22,
-91,-32,44,-43,61,56,-65,58,111,10,-21,56,-86,-56,-53,-32,-29,
25,-6,-114,24,89,-26,-14,-12,90,0,-99,0,-49,-24,3,-3,-11,




--MLP 32
/*
-157,-34,-64,-87,34,-12,-104,23,64,-26,
-98,-26,41,27,-23,14,-10,-26,-3,124,
-10,10,10,10,0,30,0,20,0,10,
-1,-30,71,-25,19,6,-67,64,39,-115,
-21,-47,73,-28,84,-54,32,-48,-46,-4,
56,106,-22,-13,-76,-149,126,-106,78,-93,
-6,4,4,12,12,2,13,3,-6,11,
57,9,-25,9,57,-47,79,14,-27,-168,
-27,-93,-128,89,60,38,-36,66,-143,144,
-48,27,-42,-16,-28,24,6,-28,-34,2,
80,-18,44,29,18,-119,15,-32,126,-145,
-15,12,10,6,-18,-24,6,23,3,20,
45,42,13,-26,-32,-2,-61,0,-42,-10,
59,14,107,-154,69,-32,-9,-74,10,4,
1,10,12,-1,3,1,2,3,13,-5,
-60,32,-78,-5,-8,-23,42,31,-18,-94,
-10,27,-16,-27,26,8,-15,32,10,9,
-8,11,2,3,21,1,2,1,11,22,
55,-14,57,-30,-52,-242,10,-71,15,133,
75,-22,18,-18,-21,120,-87,-40,-55,72,
1,11,20,9,-10,1,1,1,10,11,
-97,126,95,31,25,-70,-29,-53,-58,-170,
46,41,16,-65,-80,-18,-47,24,98,-82,
89,25,-7,-17,20,-69,-66,74,-41,29,
-49,159,-38,80,-96,17,15,54,26,-202,
79,-44,-8,-4,5,28,-63,-90,-57,29,
-46,15,37,9,-73,-35,6,35,11,69,
150,-98,-47,-49,52,18,-93,132,38,-14,
19,-102,45,-33,-68,-54,113,-22,-118,100,
-22,-2,-9,-33,17,-3,-1,-12,-7,9,
10,10,0,20,10,10,20,-10,0,-10,
-64,6,-43,-57,61,5,-9,-34,-9,102,

4697,-123,123,-44,772,1223,150,-227,402,1313,-255,198,768,-319,150,2124,297,159,1572,-666,139,2091,1133,-298,323,1276,-299,-823,634,499,118,746,

-153,10,-32,-27,-75,128,-22,-44,-12,-21,-121,16,28,-86,-22,-41,-16,-13,-86,27,-2,55,120,13,18,2,-13,51,5,-7,-22,29,-2,
123,26,-35,58,11,34,-14,-82,-81,-96,-93,-32,-18,43,-4,-50,-9,-35,98,44,-24,-29,-8,-52,-34,65,-1,6,-18,12,-16,32,-12,
134,27,-10,-28,-8,-76,-19,-61,44,-44,-103,-25,-15,-91,-9,-59,-21,-20,-38,2,-29,-113,36,32,-83,-66,1,72,-26,-32,-20,50,-8,
86,-31,-41,-24,68,73,-42,-12,80,-11,-60,-12,20,-94,-27,89,-26,-22,76,-99,-33,-52,30,14,-162,-11,-76,71,144,9,-32,1,-16,
-58,27,-5,-21,25,-17,-5,-6,-102,-23,-6,-11,-44,27,-4,-33,-4,-5,-90,26,-5,-13,6,17,-36,-17,-17,38,-16,7,5,37,4,
81,-61,-18,-70,-5,-4,-19,14,-63,-46,61,-19,14,119,-7,62,-25,-29,18,-25,-18,46,-41,34,-18,-6,-6,-50,-53,-32,-18,-14,-14,
-128,7,-14,44,-55,28,-33,-93,-68,-18,66,-28,-37,-2,-23,-1,-14,-23,93,-59,-4,-4,65,23,19,-99,-38,79,83,15,-23,61,-11,
67,47,1,-52,42,45,2,23,-111,-46,89,1,-62,-113,2,-17,14,-9,-84,-68,-9,-52,47,-79,-5,-24,-30,-43,-15,-12,1,-16,1,
-15,76,2,-12,-24,14,-18,-77,0,-5,10,-37,32,-10,-8,-4,-37,-8,10,29,-8,-84,-36,-72,18,3,59,49,23,-2,-8,-27,1,
131,49,-24,-47,-10,-105,-15,-93,-91,-30,-45,-29,42,-52,-23,87,0,-35,-88,58,-24,105,21,-7,101,-56,16,-99,-132,-33,-13,63,-4,
-14,7,6,-9,-15,-30,-33,4,19,-3,-21,17,6,-14,-3,-33,39,-14,-30,-47,6,-1,-30,-12,51,-32,-15,1,5,-12,-4,-25,5,
16,-53,3,65,-39,9,-6,28,-49,-1,-13,-5,-19,-22,-6,-9,-49,3,20,4,-17,-4,-46,-1,3,-17,41,27,-22,9,3,-21,3,
-79,15,16,-14,45,35,-13,-48,46,-41,-1,-12,-7,-69,-14,-36,14,6,-8,-45,-24,-7,-46,-14,-56,-10,-5,-45,1,-2,-14,74,4,
-47,-88,0,54,1,16,-20,9,-44,28,14,3,39,23,-29,-32,23,-19,11,48,-19,-18,40,-53,-50,42,-13,-54,-25,0,-19,-41,-7,
-26,0,-17,-111,20,-5,-17,82,38,-11,11,-35,0,-5,-26,-14,-52,-7,-9,34,-7,82,-14,73,-36,24,-60,-62,2,-14,-7,-35,-5,
*/

/*
-- MLP 64
21,1,11,11,1,1,21,11,1,1,
-6,31,21,4,-18,3,-10,28,90,-157,
-142,6,-6,-5,6,47,-20,-17,42,-24,
6,-54,169,-108,54,-35,-26,-102,36,14,
66,-18,21,10,19,27,-17,-47,-40,9,
-8,-6,-17,-1,3,-3,-24,-16,-10,28,
-2,-2,27,8,-2,8,10,20,-12,-12,
-13,22,15,-5,-3,-13,10,1,11,10,
-11,3,13,3,14,13,3,3,-8,11,
-52,27,61,-24,23,-14,1,-63,-4,-7,
-95,-2,-26,82,16,-12,-41,-59,-24,51,
-44,-7,45,11,-11,-13,-14,-16,28,7,
10,11,0,0,0,0,10,11,1,1,
10,10,10,10,0,20,11,11,-9,-9,
16,23,-61,-19,11,59,9,20,39,61,
19,-49,-17,-21,-30,-6,11,4,-18,24,
50,-104,-38,12,-110,30,32,-15,-51,65,
-71,46,14,-63,3,-15,-24,-58,57,-30,
2,55,14,-45,-9,-60,20,-50,19,-21,
-43,160,18,-11,-42,60,-38,9,-71,-153,
0,10,0,20,20,0,10,20,-10,0,
13,23,13,11,2,2,-4,13,-7,-6,
5,-75,19,-67,25,2,38,-35,33,-49,
7,18,-21,6,-27,-121,25,16,53,42,
87,20,46,-34,-62,-95,-34,-35,16,43,
0,-10,0,10,10,20,-7,11,20,11,
5,41,41,11,30,-42,5,-37,-47,-137,
69,75,0,-35,8,-33,4,-33,-88,-35,
42,-27,-40,-94,51,-14,-18,-1,-1,42,
21,8,16,-14,17,-14,7,-5,11,4,
19,29,-11,9,-1,9,-15,-1,19,0,
-62,-48,-101,10,69,51,-30,63,-105,108,
-116,16,-42,-136,51,57,-58,46,24,78,
-5,22,0,10,20,-6,-11,-13,11,-22,
-15,-11,-25,-46,-9,-6,6,28,9,15,
-10,12,-39,27,14,11,9,12,11,-21,
-6,12,1,2,2,12,13,1,20,2,
-69,-2,-42,14,0,-38,22,11,18,-42,
7,-22,-22,-12,-12,-12,-3,-12,-2,-3,
59,-12,-35,-18,67,61,-42,-57,-1,-65,
-65,-55,9,82,-40,-8,36,40,-53,-4,
-12,-8,-8,6,-9,-16,-10,1,-9,-1,
-73,-30,34,-73,32,-31,-10,2,-16,90,
2,4,-10,9,-2,8,-3,0,14,-4,
21,-25,-1,23,3,-13,-12,0,-1,-8,
-35,68,-86,-61,-37,-2,-90,19,51,25,
-36,18,-27,-41,69,1,25,24,-41,18,
-40,48,-1,-42,45,-198,11,14,61,-68,
-47,28,-42,-85,1,20,-78,179,-16,-10,
-21,4,-60,-9,-18,-4,2,1,-14,12,
-47,-22,-47,51,124,-47,26,-39,25,-85,
2,31,44,-64,-6,-31,-9,-14,35,-22,
-2,4,25,23,6,-5,5,-6,4,-3,
-78,-6,-13,38,7,58,3,27,7,-78,
-10,-8,11,79,-55,-11,61,-109,-44,46,
42,43,-6,-16,-81,-56,32,-15,125,-147,
10,9,-11,-19,21,23,-12,26,35,18,
-5,-130,11,-30,75,122,-160,14,-116,197,
3,-2,-25,-78,-5,36,-38,-87,-5,62,
0,-13,-3,-12,-15,8,-26,14,-3,-6,
-56,20,-36,12,23,48,-12,-14,27,11,
68,-21,-12,-4,14,-40,7,-14,-53,-36,
-57,42,5,-34,3,-2,-13,-49,10,-16,
22,2,12,11,-9,21,-6,11,-8,11,

142,84,1414,100,-732,357,88,144,155,613,1287,9,148,135,293,571,878,1445,565,1043,124,193,1068,281,473,140,297,653,535,198,118,489,1090,38,294,-8,157,1457,78,451,626,139,492,26,0,2241,44,2040,871,1019,481,569,204,310,562,1162,86,394,1427,223,-10,747,1067,151,


-14,-54,-51,-129,-38,-4,-4,2,7,-28,-46,-34,-14,-14,3,10,7,-88,-32,81,16,-4,-69,-10,-41,-14,17,49,-59,7,-4,-45,-51,-21,1,14,6,-69,-11,7,-42,-2,-42,-2,-29,84,26,-151,11,-43,-91,36,7,-26,55,110,-3,-26,-50,6,48,-27,-35,-14,4,
-33,-17,52,76,-28,-17,0,9,-11,19,50,-6,-12,-2,-22,-9,5,12,-42,-41,-12,-22,-8,11,9,-22,-6,-24,28,-10,-3,-91,8,-31,-3,-13,-22,-27,-1,3,-5,-5,50,-2,-5,119,-29,3,-61,-66,0,11,-1,-19,-3,45,-1,71,54,-10,9,-35,-12,-32,-2,
-22,-32,24,-68,-35,4,-1,-29,-20,-7,-2,6,-21,-2,-11,-15,0,-56,-30,-66,-22,-11,-42,10,-39,8,-24,-48,-31,-1,8,54,95,-7,-4,-8,-12,-28,-1,-1,-23,-12,-37,-17,-3,74,26,-43,95,-21,-32,2,-11,-5,-46,-27,-11,116,-59,-17,11,-47,-62,-12,-2,
-30,-71,-6,-101,-62,20,-23,-9,-21,14,-10,-11,-22,-21,-21,51,119,-44,-25,-110,-31,-12,38,41,4,-10,-33,16,17,-21,-20,50,3,-40,-3,-24,-12,36,-8,55,-1,5,-1,-45,-9,17,19,131,87,1,56,8,-14,-24,50,68,-18,124,-48,12,-39,52,-26,-20,-8,
-4,4,-7,21,4,8,-3,-1,-12,20,-58,5,-13,-4,-10,5,-25,7,-23,-28,-4,-3,-7,-3,-65,7,-26,-25,-4,-2,-24,-57,-8,0,-1,12,-3,-8,0,26,-49,9,-10,8,-8,-16,21,-25,-25,4,-21,33,8,-34,-16,18,-3,56,-42,-2,33,-23,-4,7,5,
-16,-12,-26,106,-25,9,-36,-14,-26,28,-44,0,-16,-16,-5,-10,2,22,44,21,-6,4,10,-10,3,4,-4,17,18,-33,-27,-51,-28,-27,17,19,-26,45,0,15,-18,-13,-48,-4,-3,113,-6,47,4,-34,83,-1,-15,10,-10,-21,-10,-32,-21,-1,0,14,-16,-7,7,
-9,14,-49,-54,-67,-11,21,-7,-16,2,-39,37,1,-9,23,-20,3,-40,-27,-33,1,1,-35,10,63,1,-59,22,-37,-9,0,-15,1,7,21,-12,1,-41,9,-27,-110,-2,91,-3,-9,-99,31,40,17,13,-23,28,-18,-41,-16,36,23,-41,-19,-12,51,-39,-14,1,9,
-5,68,87,-95,-37,8,-25,-23,-15,45,17,20,-5,5,7,-7,-14,-19,-39,-97,-15,-15,33,7,-56,5,-32,-60,-25,-4,-5,-69,-4,10,-18,-13,-15,14,0,31,-16,8,-23,-24,-5,34,-20,7,-50,-33,33,49,-4,35,3,68,-2,-44,-38,7,-14,-50,-14,5,6,
-24,-44,-12,10,26,-10,-4,-12,-14,-38,-19,45,6,-14,52,-11,66,-2,18,-15,-14,-14,-15,28,18,-14,-60,-8,-18,-37,-4,-25,2,18,-10,-28,-14,18,0,-53,6,-14,6,-23,7,-8,-9,-13,-17,9,-11,-35,-4,-4,18,-60,28,37,-8,10,11,-18,-13,6,8,
-14,-6,76,-34,-24,-31,-12,-4,-4,56,79,11,-14,-24,-24,-46,-87,68,31,80,-24,-23,-41,-83,-42,-24,-1,13,-82,-4,-13,-28,97,-6,-48,3,-14,20,8,-15,31,6,-68,-12,-22,84,15,-45,58,-13,-18,12,-22,62,16,-23,8,-120,-28,-14,0,-25,50,-4,3,
-14,17,-3,-26,-7,-1,-4,5,-3,-10,4,6,-4,-4,-21,-2,-14,-7,-18,10,-4,-3,-27,-7,-30,-4,-12,-21,-9,30,-4,12,-38,-2,19,-3,6,11,10,0,12,7,-12,8,-24,-28,7,-18,2,7,16,-47,-3,13,-6,0,19,-31,-28,9,27,-36,-17,-3,8,
7,58,-1,-11,22,-10,-3,-11,-1,-27,-36,-1,-3,-3,-5,20,-2,8,3,-4,-3,-13,-15,17,14,-13,6,-34,-25,-11,-13,-7,-2,-24,10,1,-3,-13,0,-11,48,28,-2,-12,7,16,-15,-16,-13,-10,-21,-48,-2,-16,14,57,5,-7,8,10,-11,-18,-2,-13,3,
-17,-27,-9,-43,-30,-12,4,-5,-6,46,40,-2,-7,3,-4,-16,-18,-18,0,-27,-7,-6,-34,9,-43,3,-28,-27,-26,-4,-17,53,-53,-4,8,-26,3,-4,10,-26,-22,9,-17,-17,-16,28,33,39,-49,-10,27,21,-15,-44,49,-14,13,13,-67,18,16,-6,-3,-7,3,
-17,5,-10,18,37,20,-7,2,-11,-2,-8,-13,-17,-17,8,-5,-12,23,23,40,-8,-17,-5,19,7,-18,36,34,6,3,-7,-26,-34,-7,8,-30,-27,-19,-20,74,-42,10,-24,-8,-15,-23,-63,-46,-28,8,-31,36,-17,-12,1,16,-24,-3,-16,-21,-3,25,25,13,5,
-6,-94,-27,-35,12,19,14,-17,5,-7,17,-27,4,14,-47,11,-70,18,11,-9,4,4,-22,-27,-6,-16,44,36,26,24,-16,-8,-16,2,0,9,3,-21,10,46,-2,16,-4,4,26,14,-14,-6,-4,10,1,-29,13,15,4,-42,-22,-45,26,-10,-29,45,-2,-16,33,
*/


others => 0
    );
    
begin

process(all)  --data memory
begin
if rising_edge(clk) then
    if READ_RAM = '1' then --read data from RAM memory
        DATA_RAM_OUT <= std_logic_vector(to_signed(RAM_DATA(to_integer(unsigned(ADDRESS_DATA))),data)) after 10 ns;
    elsif WRITE_RAM = '1' then --write data to RAM memory
        RAM_DATA(to_integer(unsigned(ADDRESS_DATA))) <= to_integer(signed(DATA_RAM_IN));
    elsif WRITE_RESET = '1' then
        RAM_DATA(to_integer(unsigned(RESET_ADDRESS))) <= to_integer(signed(RESET_DATA)); 
    end if;
end if;
end process;
end Behavioral;

