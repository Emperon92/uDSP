library IEEE;

use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.std_logic_unsigned.all;

package walltree_func is
    function mul_func ( 
        OP1_mul: in std_logic_vector(15 downto 0 );
        OP2_mul: in std_logic_vector(15 downto 0 ))
        return std_logic_vector;
end package walltree_func;

package body walltree_func is

 function mul_func (
    OP1_mul: in std_logic_vector(15 downto 0 );
    OP2_mul: in std_logic_vector(15 downto 0 ))
    return std_logic_vector is
    
        variable pp0 : std_logic_vector(15 downto 0 );
        variable  pp1 : std_logic_vector(15 downto 0 );
        variable  pp2 : std_logic_vector(15 downto 0 );
        variable  pp3 : std_logic_vector(15 downto 0 );
        variable  pp4 : std_logic_vector(15 downto 0 );
        variable  pp5 : std_logic_vector(15 downto 0 );
        variable  pp6 : std_logic_vector(15 downto 0 );
        variable  pp7 : std_logic_vector(15 downto 0 );
        variable  pp8 : std_logic_vector(15 downto 0 );
        variable  pp9 : std_logic_vector(15 downto 0 );
        variable  pp10 : std_logic_vector(15 downto 0 );
        variable  pp11 : std_logic_vector(15 downto 0 );
        variable  pp12 : std_logic_vector(15 downto 0 );
        variable  pp13 : std_logic_vector(15 downto 0 );
        variable  pp14 : std_logic_vector(15 downto 0 );
        variable  pp15 : std_logic_vector(15 downto 0 );
        
        -- internal signals

        -- layer : 1
        
        -- csa : 0
        variable sigCSA_sum_0 : std_logic_vector (17 downto 0);
        variable sigCSA_cry_0 : std_logic_vector (17 downto 0);
        -- csa : 1
        variable sigCSA_sum_1 : std_logic_vector (17 downto 0);
        variable sigCSA_cry_1 : std_logic_vector (17 downto 0);
        -- csa : 2
        variable sigCSA_sum_2 : std_logic_vector (17 downto 0);
        variable sigCSA_cry_2 : std_logic_vector (17 downto 0);
        -- csa : 3
        variable sigCSA_sum_3 : std_logic_vector (17 downto 0);
        variable sigCSA_cry_3 : std_logic_vector (17 downto 0);
        -- csa : 4
        variable sigCSA_sum_4 : std_logic_vector (17 downto 0);
        variable sigCSA_cry_4 : std_logic_vector (17 downto 0);
        
        -- layer : 2
        
        -- csa : 5
        variable sigCSA_sum_5 : std_logic_vector (20 downto 0);
        variable sigCSA_cry_5 : std_logic_vector (20 downto 0);
        -- csa : 6
        variable sigCSA_sum_6 : std_logic_vector (20 downto 0);
        variable sigCSA_cry_6 : std_logic_vector (20 downto 0);
        -- csa : 7
        variable sigCSA_sum_7 : std_logic_vector (20 downto 0);
        variable sigCSA_cry_7 : std_logic_vector (20 downto 0);
        
        -- layer : 3
        
        -- csa : 8
        variable sigCSA_sum_8 : std_logic_vector (24 downto 0);
        variable sigCSA_cry_8 : std_logic_vector (24 downto 0);
        -- csa : 9
        variable sigCSA_sum_9 : std_logic_vector (25 downto 0);
        variable sigCSA_cry_9 : std_logic_vector (25 downto 0);
        
        -- layer : 4
        
        -- csa : 10
        variable sigCSA_sum_10 : std_logic_vector (30 downto 0);
        variable sigCSA_cry_10 : std_logic_vector (30 downto 0);
        -- csa : 11
        variable sigCSA_sum_11 : std_logic_vector (30 downto 0);
        variable sigCSA_cry_11 : std_logic_vector (30 downto 0);
        
        -- layer : 5
        
        -- csa : 12
        variable sigCSA_sum_12 : std_logic_vector (32 downto 0);
        variable sigCSA_cry_12 : std_logic_vector (32 downto 0);
        
        -- layer : 6
        
        -- csa : 13
        variable sigCSA_sum_13 : std_logic_vector (32 downto 0);
        variable sigCSA_cry_13 : std_logic_vector (32 downto 0);
        --sigCSA_sum_13
        --sigCSA_cry_13
        -- all csa structures generated
        -- carry variable for the final RCA
        
        variable carry_rca : std_logic_vector(31 downto 0 );
        
        variable result_int : std_logic_vector(32 downto 0 );
        
        begin 
        
        --walltree_mul

        pp0(0) := OP1_mul(0) and OP2_mul(0);
        pp0(1) := OP1_mul(0) and OP2_mul(1);
        pp0(2) := OP1_mul(0) and OP2_mul(2);
        pp0(3) := OP1_mul(0) and OP2_mul(3);
        pp0(4) := OP1_mul(0) and OP2_mul(4);
        pp0(5) := OP1_mul(0) and OP2_mul(5);
        pp0(6) := OP1_mul(0) and OP2_mul(6);
        pp0(7) := OP1_mul(0) and OP2_mul(7);
        pp0(8) := OP1_mul(0) and OP2_mul(8);
        pp0(9) := OP1_mul(0) and OP2_mul(9);
        pp0(10) := OP1_mul(0) and OP2_mul(10);
        pp0(11) := OP1_mul(0) and OP2_mul(11);
        pp0(12) := OP1_mul(0) and OP2_mul(12);
        pp0(13) := OP1_mul(0) and OP2_mul(13);
        pp0(14) := OP1_mul(0) and OP2_mul(14);
        pp0(15) := OP1_mul(0) and OP2_mul(15);
        pp1(0) := OP1_mul(1) and OP2_mul(0);
        pp1(1) := OP1_mul(1) and OP2_mul(1);
        pp1(2) := OP1_mul(1) and OP2_mul(2);
        pp1(3) := OP1_mul(1) and OP2_mul(3);
        pp1(4) := OP1_mul(1) and OP2_mul(4);
        pp1(5) := OP1_mul(1) and OP2_mul(5);
        pp1(6) := OP1_mul(1) and OP2_mul(6);
        pp1(7) := OP1_mul(1) and OP2_mul(7);
        pp1(8) := OP1_mul(1) and OP2_mul(8);
        pp1(9) := OP1_mul(1) and OP2_mul(9);
        pp1(10) := OP1_mul(1) and OP2_mul(10);
        pp1(11) := OP1_mul(1) and OP2_mul(11);
        pp1(12) := OP1_mul(1) and OP2_mul(12);
        pp1(13) := OP1_mul(1) and OP2_mul(13);
        pp1(14) := OP1_mul(1) and OP2_mul(14);
        pp1(15) := OP1_mul(1) and OP2_mul(15);
        pp2(0) := OP1_mul(2) and OP2_mul(0);
        pp2(1) := OP1_mul(2) and OP2_mul(1);
        pp2(2) := OP1_mul(2) and OP2_mul(2);
        pp2(3) := OP1_mul(2) and OP2_mul(3);
        pp2(4) := OP1_mul(2) and OP2_mul(4);
        pp2(5) := OP1_mul(2) and OP2_mul(5);
        pp2(6) := OP1_mul(2) and OP2_mul(6);
        pp2(7) := OP1_mul(2) and OP2_mul(7);
        pp2(8) := OP1_mul(2) and OP2_mul(8);
        pp2(9) := OP1_mul(2) and OP2_mul(9);
        pp2(10) := OP1_mul(2) and OP2_mul(10);
        pp2(11) := OP1_mul(2) and OP2_mul(11);
        pp2(12) := OP1_mul(2) and OP2_mul(12);
        pp2(13) := OP1_mul(2) and OP2_mul(13);
        pp2(14) := OP1_mul(2) and OP2_mul(14);
        pp2(15) := OP1_mul(2) and OP2_mul(15);
        pp3(0) := OP1_mul(3) and OP2_mul(0);
        pp3(1) := OP1_mul(3) and OP2_mul(1);
        pp3(2) := OP1_mul(3) and OP2_mul(2);
        pp3(3) := OP1_mul(3) and OP2_mul(3);
        pp3(4) := OP1_mul(3) and OP2_mul(4);
        pp3(5) := OP1_mul(3) and OP2_mul(5);
        pp3(6) := OP1_mul(3) and OP2_mul(6);
        pp3(7) := OP1_mul(3) and OP2_mul(7);
        pp3(8) := OP1_mul(3) and OP2_mul(8);
        pp3(9) := OP1_mul(3) and OP2_mul(9);
        pp3(10) := OP1_mul(3) and OP2_mul(10);
        pp3(11) := OP1_mul(3) and OP2_mul(11);
        pp3(12) := OP1_mul(3) and OP2_mul(12);
        pp3(13) := OP1_mul(3) and OP2_mul(13);
        pp3(14) := OP1_mul(3) and OP2_mul(14);
        pp3(15) := OP1_mul(3) and OP2_mul(15);
        pp4(0) := OP1_mul(4) and OP2_mul(0);
        pp4(1) := OP1_mul(4) and OP2_mul(1);
        pp4(2) := OP1_mul(4) and OP2_mul(2);
        pp4(3) := OP1_mul(4) and OP2_mul(3);
        pp4(4) := OP1_mul(4) and OP2_mul(4);
        pp4(5) := OP1_mul(4) and OP2_mul(5);
        pp4(6) := OP1_mul(4) and OP2_mul(6);
        pp4(7) := OP1_mul(4) and OP2_mul(7);
        pp4(8) := OP1_mul(4) and OP2_mul(8);
        pp4(9) := OP1_mul(4) and OP2_mul(9);
        pp4(10) := OP1_mul(4) and OP2_mul(10);
        pp4(11) := OP1_mul(4) and OP2_mul(11);
        pp4(12) := OP1_mul(4) and OP2_mul(12);
        pp4(13) := OP1_mul(4) and OP2_mul(13);
        pp4(14) := OP1_mul(4) and OP2_mul(14);
        pp4(15) := OP1_mul(4) and OP2_mul(15);
        pp5(0) := OP1_mul(5) and OP2_mul(0);
        pp5(1) := OP1_mul(5) and OP2_mul(1);
        pp5(2) := OP1_mul(5) and OP2_mul(2);
        pp5(3) := OP1_mul(5) and OP2_mul(3);
        pp5(4) := OP1_mul(5) and OP2_mul(4);
        pp5(5) := OP1_mul(5) and OP2_mul(5);
        pp5(6) := OP1_mul(5) and OP2_mul(6);
        pp5(7) := OP1_mul(5) and OP2_mul(7);
        pp5(8) := OP1_mul(5) and OP2_mul(8);
        pp5(9) := OP1_mul(5) and OP2_mul(9);
        pp5(10) := OP1_mul(5) and OP2_mul(10);
        pp5(11) := OP1_mul(5) and OP2_mul(11);
        pp5(12) := OP1_mul(5) and OP2_mul(12);
        pp5(13) := OP1_mul(5) and OP2_mul(13);
        pp5(14) := OP1_mul(5) and OP2_mul(14);
        pp5(15) := OP1_mul(5) and OP2_mul(15);
        pp6(0) := OP1_mul(6) and OP2_mul(0);
        pp6(1) := OP1_mul(6) and OP2_mul(1);
        pp6(2) := OP1_mul(6) and OP2_mul(2);
        pp6(3) := OP1_mul(6) and OP2_mul(3);
        pp6(4) := OP1_mul(6) and OP2_mul(4);
        pp6(5) := OP1_mul(6) and OP2_mul(5);
        pp6(6) := OP1_mul(6) and OP2_mul(6);
        pp6(7) := OP1_mul(6) and OP2_mul(7);
        pp6(8) := OP1_mul(6) and OP2_mul(8);
        pp6(9) := OP1_mul(6) and OP2_mul(9);
        pp6(10) := OP1_mul(6) and OP2_mul(10);
        pp6(11) := OP1_mul(6) and OP2_mul(11);
        pp6(12) := OP1_mul(6) and OP2_mul(12);
        pp6(13) := OP1_mul(6) and OP2_mul(13);
        pp6(14) := OP1_mul(6) and OP2_mul(14);
        pp6(15) := OP1_mul(6) and OP2_mul(15);
        pp7(0) := OP1_mul(7) and OP2_mul(0);
        pp7(1) := OP1_mul(7) and OP2_mul(1);
        pp7(2) := OP1_mul(7) and OP2_mul(2);
        pp7(3) := OP1_mul(7) and OP2_mul(3);
        pp7(4) := OP1_mul(7) and OP2_mul(4);
        pp7(5) := OP1_mul(7) and OP2_mul(5);
        pp7(6) := OP1_mul(7) and OP2_mul(6);
        pp7(7) := OP1_mul(7) and OP2_mul(7);
        pp7(8) := OP1_mul(7) and OP2_mul(8);
        pp7(9) := OP1_mul(7) and OP2_mul(9);
        pp7(10) := OP1_mul(7) and OP2_mul(10);
        pp7(11) := OP1_mul(7) and OP2_mul(11);
        pp7(12) := OP1_mul(7) and OP2_mul(12);
        pp7(13) := OP1_mul(7) and OP2_mul(13);
        pp7(14) := OP1_mul(7) and OP2_mul(14);
        pp7(15) := OP1_mul(7) and OP2_mul(15);
        pp8(0) := OP1_mul(8) and OP2_mul(0);
        pp8(1) := OP1_mul(8) and OP2_mul(1);
        pp8(2) := OP1_mul(8) and OP2_mul(2);
        pp8(3) := OP1_mul(8) and OP2_mul(3);
        pp8(4) := OP1_mul(8) and OP2_mul(4);
        pp8(5) := OP1_mul(8) and OP2_mul(5);
        pp8(6) := OP1_mul(8) and OP2_mul(6);
        pp8(7) := OP1_mul(8) and OP2_mul(7);
        pp8(8) := OP1_mul(8) and OP2_mul(8);
        pp8(9) := OP1_mul(8) and OP2_mul(9);
        pp8(10) := OP1_mul(8) and OP2_mul(10);
        pp8(11) := OP1_mul(8) and OP2_mul(11);
        pp8(12) := OP1_mul(8) and OP2_mul(12);
        pp8(13) := OP1_mul(8) and OP2_mul(13);
        pp8(14) := OP1_mul(8) and OP2_mul(14);
        pp8(15) := OP1_mul(8) and OP2_mul(15);
        pp9(0) := OP1_mul(9) and OP2_mul(0);
        pp9(1) := OP1_mul(9) and OP2_mul(1);
        pp9(2) := OP1_mul(9) and OP2_mul(2);
        pp9(3) := OP1_mul(9) and OP2_mul(3);
        pp9(4) := OP1_mul(9) and OP2_mul(4);
        pp9(5) := OP1_mul(9) and OP2_mul(5);
        pp9(6) := OP1_mul(9) and OP2_mul(6);
        pp9(7) := OP1_mul(9) and OP2_mul(7);
        pp9(8) := OP1_mul(9) and OP2_mul(8);
        pp9(9) := OP1_mul(9) and OP2_mul(9);
        pp9(10) := OP1_mul(9) and OP2_mul(10);
        pp9(11) := OP1_mul(9) and OP2_mul(11);
        pp9(12) := OP1_mul(9) and OP2_mul(12);
        pp9(13) := OP1_mul(9) and OP2_mul(13);
        pp9(14) := OP1_mul(9) and OP2_mul(14);
        pp9(15) := OP1_mul(9) and OP2_mul(15);
        pp10(0) := OP1_mul(10) and OP2_mul(0);
        pp10(1) := OP1_mul(10) and OP2_mul(1);
        pp10(2) := OP1_mul(10) and OP2_mul(2);
        pp10(3) := OP1_mul(10) and OP2_mul(3);
        pp10(4) := OP1_mul(10) and OP2_mul(4);
        pp10(5) := OP1_mul(10) and OP2_mul(5);
        pp10(6) := OP1_mul(10) and OP2_mul(6);
        pp10(7) := OP1_mul(10) and OP2_mul(7);
        pp10(8) := OP1_mul(10) and OP2_mul(8);
        pp10(9) := OP1_mul(10) and OP2_mul(9);
        pp10(10) := OP1_mul(10) and OP2_mul(10);
        pp10(11) := OP1_mul(10) and OP2_mul(11);
        pp10(12) := OP1_mul(10) and OP2_mul(12);
        pp10(13) := OP1_mul(10) and OP2_mul(13);
        pp10(14) := OP1_mul(10) and OP2_mul(14);
        pp10(15) := OP1_mul(10) and OP2_mul(15);
        pp11(0) := OP1_mul(11) and OP2_mul(0);
        pp11(1) := OP1_mul(11) and OP2_mul(1);
        pp11(2) := OP1_mul(11) and OP2_mul(2);
        pp11(3) := OP1_mul(11) and OP2_mul(3);
        pp11(4) := OP1_mul(11) and OP2_mul(4);
        pp11(5) := OP1_mul(11) and OP2_mul(5);
        pp11(6) := OP1_mul(11) and OP2_mul(6);
        pp11(7) := OP1_mul(11) and OP2_mul(7);
        pp11(8) := OP1_mul(11) and OP2_mul(8);
        pp11(9) := OP1_mul(11) and OP2_mul(9);
        pp11(10) := OP1_mul(11) and OP2_mul(10);
        pp11(11) := OP1_mul(11) and OP2_mul(11);
        pp11(12) := OP1_mul(11) and OP2_mul(12);
        pp11(13) := OP1_mul(11) and OP2_mul(13);
        pp11(14) := OP1_mul(11) and OP2_mul(14);
        pp11(15) := OP1_mul(11) and OP2_mul(15);
        pp12(0) := OP1_mul(12) and OP2_mul(0);
        pp12(1) := OP1_mul(12) and OP2_mul(1);
        pp12(2) := OP1_mul(12) and OP2_mul(2);
        pp12(3) := OP1_mul(12) and OP2_mul(3);
        pp12(4) := OP1_mul(12) and OP2_mul(4);
        pp12(5) := OP1_mul(12) and OP2_mul(5);
        pp12(6) := OP1_mul(12) and OP2_mul(6);
        pp12(7) := OP1_mul(12) and OP2_mul(7);
        pp12(8) := OP1_mul(12) and OP2_mul(8);
        pp12(9) := OP1_mul(12) and OP2_mul(9);
        pp12(10) := OP1_mul(12) and OP2_mul(10);
        pp12(11) := OP1_mul(12) and OP2_mul(11);
        pp12(12) := OP1_mul(12) and OP2_mul(12);
        pp12(13) := OP1_mul(12) and OP2_mul(13);
        pp12(14) := OP1_mul(12) and OP2_mul(14);
        pp12(15) := OP1_mul(12) and OP2_mul(15);
        pp13(0) := OP1_mul(13) and OP2_mul(0);
        pp13(1) := OP1_mul(13) and OP2_mul(1);
        pp13(2) := OP1_mul(13) and OP2_mul(2);
        pp13(3) := OP1_mul(13) and OP2_mul(3);
        pp13(4) := OP1_mul(13) and OP2_mul(4);
        pp13(5) := OP1_mul(13) and OP2_mul(5);
        pp13(6) := OP1_mul(13) and OP2_mul(6);
        pp13(7) := OP1_mul(13) and OP2_mul(7);
        pp13(8) := OP1_mul(13) and OP2_mul(8);
        pp13(9) := OP1_mul(13) and OP2_mul(9);
        pp13(10) := OP1_mul(13) and OP2_mul(10);
        pp13(11) := OP1_mul(13) and OP2_mul(11);
        pp13(12) := OP1_mul(13) and OP2_mul(12);
        pp13(13) := OP1_mul(13) and OP2_mul(13);
        pp13(14) := OP1_mul(13) and OP2_mul(14);
        pp13(15) := OP1_mul(13) and OP2_mul(15);
        pp14(0) := OP1_mul(14) and OP2_mul(0);
        pp14(1) := OP1_mul(14) and OP2_mul(1);
        pp14(2) := OP1_mul(14) and OP2_mul(2);
        pp14(3) := OP1_mul(14) and OP2_mul(3);
        pp14(4) := OP1_mul(14) and OP2_mul(4);
        pp14(5) := OP1_mul(14) and OP2_mul(5);
        pp14(6) := OP1_mul(14) and OP2_mul(6);
        pp14(7) := OP1_mul(14) and OP2_mul(7);
        pp14(8) := OP1_mul(14) and OP2_mul(8);
        pp14(9) := OP1_mul(14) and OP2_mul(9);
        pp14(10) := OP1_mul(14) and OP2_mul(10);
        pp14(11) := OP1_mul(14) and OP2_mul(11);
        pp14(12) := OP1_mul(14) and OP2_mul(12);
        pp14(13) := OP1_mul(14) and OP2_mul(13);
        pp14(14) := OP1_mul(14) and OP2_mul(14);
        pp14(15) := OP1_mul(14) and OP2_mul(15);
        pp15(0) := OP1_mul(15) and OP2_mul(0);
        pp15(1) := OP1_mul(15) and OP2_mul(1);
        pp15(2) := OP1_mul(15) and OP2_mul(2);
        pp15(3) := OP1_mul(15) and OP2_mul(3);
        pp15(4) := OP1_mul(15) and OP2_mul(4);
        pp15(5) := OP1_mul(15) and OP2_mul(5);
        pp15(6) := OP1_mul(15) and OP2_mul(6);
        pp15(7) := OP1_mul(15) and OP2_mul(7);
        pp15(8) := OP1_mul(15) and OP2_mul(8);
        pp15(9) := OP1_mul(15) and OP2_mul(9);
        pp15(10) := OP1_mul(15) and OP2_mul(10);
        pp15(11) := OP1_mul(15) and OP2_mul(11);
        pp15(12) := OP1_mul(15) and OP2_mul(12);
        pp15(13) := OP1_mul(15) and OP2_mul(13);
        pp15(14) := OP1_mul(15) and OP2_mul(14);
        pp15(15) := OP1_mul(15) and OP2_mul(15);
-- ******************
-- csa : 0
-- generating sigCSA_sum_0 and sigCSA_cry_0

        sigCSA_sum_0(0) := pp0(0) xor '0' xor '0' ;
        sigCSA_cry_0(0) := ( pp0(0) and '0' ) or ( '0' and ( pp0(0) xor '0' )) ;
        sigCSA_sum_0(1) := pp0(1) xor pp1(0) xor '0' ;
        sigCSA_cry_0(1) := ( pp0(1) and pp1(0) ) or ( '0' and ( pp0(1) xor pp1(0) )) ;
        sigCSA_sum_0(2) := pp0(2) xor pp1(1) xor pp2(0) ;
        sigCSA_cry_0(2) := ( pp0(2) and pp1(1) ) or ( pp2(0) and ( pp0(2) xor pp1(1) )) ;
        sigCSA_sum_0(3) := pp0(3) xor pp1(2) xor pp2(1) ;
        sigCSA_cry_0(3) := ( pp0(3) and pp1(2) ) or ( pp2(1) and ( pp0(3) xor pp1(2) )) ;
        sigCSA_sum_0(4) := pp0(4) xor pp1(3) xor pp2(2) ;
        sigCSA_cry_0(4) := ( pp0(4) and pp1(3) ) or ( pp2(2) and ( pp0(4) xor pp1(3) )) ;
        sigCSA_sum_0(5) := pp0(5) xor pp1(4) xor pp2(3) ;
        sigCSA_cry_0(5) := ( pp0(5) and pp1(4) ) or ( pp2(3) and ( pp0(5) xor pp1(4) )) ;
        sigCSA_sum_0(6) := pp0(6) xor pp1(5) xor pp2(4) ;
        sigCSA_cry_0(6) := ( pp0(6) and pp1(5) ) or ( pp2(4) and ( pp0(6) xor pp1(5) )) ;
        sigCSA_sum_0(7) := pp0(7) xor pp1(6) xor pp2(5) ;
        sigCSA_cry_0(7) := ( pp0(7) and pp1(6) ) or ( pp2(5) and ( pp0(7) xor pp1(6) )) ;
        sigCSA_sum_0(8) := pp0(8) xor pp1(7) xor pp2(6) ;
        sigCSA_cry_0(8) := ( pp0(8) and pp1(7) ) or ( pp2(6) and ( pp0(8) xor pp1(7) )) ;
        sigCSA_sum_0(9) := pp0(9) xor pp1(8) xor pp2(7) ;
        sigCSA_cry_0(9) := ( pp0(9) and pp1(8) ) or ( pp2(7) and ( pp0(9) xor pp1(8) )) ;
        sigCSA_sum_0(10) := pp0(10) xor pp1(9) xor pp2(8) ;
        sigCSA_cry_0(10) := ( pp0(10) and pp1(9) ) or ( pp2(8) and ( pp0(10) xor pp1(9) )) ;
        sigCSA_sum_0(11) := pp0(11) xor pp1(10) xor pp2(9) ;
        sigCSA_cry_0(11) := ( pp0(11) and pp1(10) ) or ( pp2(9) and ( pp0(11) xor pp1(10) )) ;
        sigCSA_sum_0(12) := pp0(12) xor pp1(11) xor pp2(10) ;
        sigCSA_cry_0(12) := ( pp0(12) and pp1(11) ) or ( pp2(10) and ( pp0(12) xor pp1(11) )) ;
        sigCSA_sum_0(13) := pp0(13) xor pp1(12) xor pp2(11) ;
        sigCSA_cry_0(13) := ( pp0(13) and pp1(12) ) or ( pp2(11) and ( pp0(13) xor pp1(12) )) ;
        sigCSA_sum_0(14) := pp0(14) xor pp1(13) xor pp2(12) ;
        sigCSA_cry_0(14) := ( pp0(14) and pp1(13) ) or ( pp2(12) and ( pp0(14) xor pp1(13) )) ;
        sigCSA_sum_0(15) := pp0(15) xor pp1(14) xor pp2(13) ;
        sigCSA_cry_0(15) := ( pp0(15) and pp1(14) ) or ( pp2(13) and ( pp0(15) xor pp1(14) )) ;
        sigCSA_sum_0(16) := '0' xor pp1(15) xor pp2(14) ;
        sigCSA_cry_0(16) := ( '0' and pp1(15) ) or ( pp2(14) and ( '0' xor pp1(15) )) ;
        sigCSA_sum_0(17) := '0' xor '0' xor pp2(15) ;
        sigCSA_cry_0(17) := ( '0' and '0' ) or ( pp2(15) and ( '0' xor '0' )) ;
-- csa : 1
-- generating sigCSA_sum_1 and sigCSA_cry_1

        sigCSA_sum_1(0) := pp3(0) xor '0' xor '0' ;
        sigCSA_cry_1(0) := ( pp3(0) and '0' ) or ( '0' and ( pp3(0) xor '0' )) ;
        sigCSA_sum_1(1) := pp3(1) xor pp4(0) xor '0' ;
        sigCSA_cry_1(1) := ( pp3(1) and pp4(0) ) or ( '0' and ( pp3(1) xor pp4(0) )) ;
        sigCSA_sum_1(2) := pp3(2) xor pp4(1) xor pp5(0) ;
        sigCSA_cry_1(2) := ( pp3(2) and pp4(1) ) or ( pp5(0) and ( pp3(2) xor pp4(1) )) ;
        sigCSA_sum_1(3) := pp3(3) xor pp4(2) xor pp5(1) ;
        sigCSA_cry_1(3) := ( pp3(3) and pp4(2) ) or ( pp5(1) and ( pp3(3) xor pp4(2) )) ;
        sigCSA_sum_1(4) := pp3(4) xor pp4(3) xor pp5(2) ;
        sigCSA_cry_1(4) := ( pp3(4) and pp4(3) ) or ( pp5(2) and ( pp3(4) xor pp4(3) )) ;
        sigCSA_sum_1(5) := pp3(5) xor pp4(4) xor pp5(3) ;
        sigCSA_cry_1(5) := ( pp3(5) and pp4(4) ) or ( pp5(3) and ( pp3(5) xor pp4(4) )) ;
        sigCSA_sum_1(6) := pp3(6) xor pp4(5) xor pp5(4) ;
        sigCSA_cry_1(6) := ( pp3(6) and pp4(5) ) or ( pp5(4) and ( pp3(6) xor pp4(5) )) ;
        sigCSA_sum_1(7) := pp3(7) xor pp4(6) xor pp5(5) ;
        sigCSA_cry_1(7) := ( pp3(7) and pp4(6) ) or ( pp5(5) and ( pp3(7) xor pp4(6) )) ;
        sigCSA_sum_1(8) := pp3(8) xor pp4(7) xor pp5(6) ;
        sigCSA_cry_1(8) := ( pp3(8) and pp4(7) ) or ( pp5(6) and ( pp3(8) xor pp4(7) )) ;
        sigCSA_sum_1(9) := pp3(9) xor pp4(8) xor pp5(7) ;
        sigCSA_cry_1(9) := ( pp3(9) and pp4(8) ) or ( pp5(7) and ( pp3(9) xor pp4(8) )) ;
        sigCSA_sum_1(10) := pp3(10) xor pp4(9) xor pp5(8) ;
        sigCSA_cry_1(10) := ( pp3(10) and pp4(9) ) or ( pp5(8) and ( pp3(10) xor pp4(9) )) ;
        sigCSA_sum_1(11) := pp3(11) xor pp4(10) xor pp5(9) ;
        sigCSA_cry_1(11) := ( pp3(11) and pp4(10) ) or ( pp5(9) and ( pp3(11) xor pp4(10) )) ;
        sigCSA_sum_1(12) := pp3(12) xor pp4(11) xor pp5(10) ;
        sigCSA_cry_1(12) := ( pp3(12) and pp4(11) ) or ( pp5(10) and ( pp3(12) xor pp4(11) )) ;
        sigCSA_sum_1(13) := pp3(13) xor pp4(12) xor pp5(11) ;
        sigCSA_cry_1(13) := ( pp3(13) and pp4(12) ) or ( pp5(11) and ( pp3(13) xor pp4(12) )) ;
        sigCSA_sum_1(14) := pp3(14) xor pp4(13) xor pp5(12) ;
        sigCSA_cry_1(14) := ( pp3(14) and pp4(13) ) or ( pp5(12) and ( pp3(14) xor pp4(13) )) ;
        sigCSA_sum_1(15) := pp3(15) xor pp4(14) xor pp5(13) ;
        sigCSA_cry_1(15) := ( pp3(15) and pp4(14) ) or ( pp5(13) and ( pp3(15) xor pp4(14) )) ;
        sigCSA_sum_1(16) := '0' xor pp4(15) xor pp5(14) ;
        sigCSA_cry_1(16) := ( '0' and pp4(15) ) or ( pp5(14) and ( '0' xor pp4(15) )) ;
        sigCSA_sum_1(17) := '0' xor '0' xor pp5(15) ;
        sigCSA_cry_1(17) := ( '0' and '0' ) or ( pp5(15) and ( '0' xor '0' )) ;
-- csa : 2
-- generating sigCSA_sum_2 and sigCSA_cry_2

        sigCSA_sum_2(0) := pp6(0) xor '0' xor '0' ;
        sigCSA_cry_2(0) := ( pp6(0) and '0' ) or ( '0' and ( pp6(0) xor '0' )) ;
        sigCSA_sum_2(1) := pp6(1) xor pp7(0) xor '0' ;
        sigCSA_cry_2(1) := ( pp6(1) and pp7(0) ) or ( '0' and ( pp6(1) xor pp7(0) )) ;
        sigCSA_sum_2(2) := pp6(2) xor pp7(1) xor pp8(0) ;
        sigCSA_cry_2(2) := ( pp6(2) and pp7(1) ) or ( pp8(0) and ( pp6(2) xor pp7(1) )) ;
        sigCSA_sum_2(3) := pp6(3) xor pp7(2) xor pp8(1) ;
        sigCSA_cry_2(3) := ( pp6(3) and pp7(2) ) or ( pp8(1) and ( pp6(3) xor pp7(2) )) ;
        sigCSA_sum_2(4) := pp6(4) xor pp7(3) xor pp8(2) ;
        sigCSA_cry_2(4) := ( pp6(4) and pp7(3) ) or ( pp8(2) and ( pp6(4) xor pp7(3) )) ;
        sigCSA_sum_2(5) := pp6(5) xor pp7(4) xor pp8(3) ;
        sigCSA_cry_2(5) := ( pp6(5) and pp7(4) ) or ( pp8(3) and ( pp6(5) xor pp7(4) )) ;
        sigCSA_sum_2(6) := pp6(6) xor pp7(5) xor pp8(4) ;
        sigCSA_cry_2(6) := ( pp6(6) and pp7(5) ) or ( pp8(4) and ( pp6(6) xor pp7(5) )) ;
        sigCSA_sum_2(7) := pp6(7) xor pp7(6) xor pp8(5) ;
        sigCSA_cry_2(7) := ( pp6(7) and pp7(6) ) or ( pp8(5) and ( pp6(7) xor pp7(6) )) ;
        sigCSA_sum_2(8) := pp6(8) xor pp7(7) xor pp8(6) ;
        sigCSA_cry_2(8) := ( pp6(8) and pp7(7) ) or ( pp8(6) and ( pp6(8) xor pp7(7) )) ;
        sigCSA_sum_2(9) := pp6(9) xor pp7(8) xor pp8(7) ;
        sigCSA_cry_2(9) := ( pp6(9) and pp7(8) ) or ( pp8(7) and ( pp6(9) xor pp7(8) )) ;
        sigCSA_sum_2(10) := pp6(10) xor pp7(9) xor pp8(8) ;
        sigCSA_cry_2(10) := ( pp6(10) and pp7(9) ) or ( pp8(8) and ( pp6(10) xor pp7(9) )) ;
        sigCSA_sum_2(11) := pp6(11) xor pp7(10) xor pp8(9) ;
        sigCSA_cry_2(11) := ( pp6(11) and pp7(10) ) or ( pp8(9) and ( pp6(11) xor pp7(10) )) ;
        sigCSA_sum_2(12) := pp6(12) xor pp7(11) xor pp8(10) ;
        sigCSA_cry_2(12) := ( pp6(12) and pp7(11) ) or ( pp8(10) and ( pp6(12) xor pp7(11) )) ;
        sigCSA_sum_2(13) := pp6(13) xor pp7(12) xor pp8(11) ;
        sigCSA_cry_2(13) := ( pp6(13) and pp7(12) ) or ( pp8(11) and ( pp6(13) xor pp7(12) )) ;
        sigCSA_sum_2(14) := pp6(14) xor pp7(13) xor pp8(12) ;
        sigCSA_cry_2(14) := ( pp6(14) and pp7(13) ) or ( pp8(12) and ( pp6(14) xor pp7(13) )) ;
        sigCSA_sum_2(15) := pp6(15) xor pp7(14) xor pp8(13) ;
        sigCSA_cry_2(15) := ( pp6(15) and pp7(14) ) or ( pp8(13) and ( pp6(15) xor pp7(14) )) ;
        sigCSA_sum_2(16) := '0' xor pp7(15) xor pp8(14) ;
        sigCSA_cry_2(16) := ( '0' and pp7(15) ) or ( pp8(14) and ( '0' xor pp7(15) )) ;
        sigCSA_sum_2(17) := '0' xor '0' xor pp8(15) ;
        sigCSA_cry_2(17) := ( '0' and '0' ) or ( pp8(15) and ( '0' xor '0' )) ;
-- csa : 3
-- generating sigCSA_sum_3 and sigCSA_cry_3

        sigCSA_sum_3(0) := pp9(0) xor '0' xor '0' ;
        sigCSA_cry_3(0) := ( pp9(0) and '0' ) or ( '0' and ( pp9(0) xor '0' )) ;
        sigCSA_sum_3(1) := pp9(1) xor pp10(0) xor '0' ;
        sigCSA_cry_3(1) := ( pp9(1) and pp10(0) ) or ( '0' and ( pp9(1) xor pp10(0) )) ;
        sigCSA_sum_3(2) := pp9(2) xor pp10(1) xor pp11(0) ;
        sigCSA_cry_3(2) := ( pp9(2) and pp10(1) ) or ( pp11(0) and ( pp9(2) xor pp10(1) )) ;
        sigCSA_sum_3(3) := pp9(3) xor pp10(2) xor pp11(1) ;
        sigCSA_cry_3(3) := ( pp9(3) and pp10(2) ) or ( pp11(1) and ( pp9(3) xor pp10(2) )) ;
        sigCSA_sum_3(4) := pp9(4) xor pp10(3) xor pp11(2) ;
        sigCSA_cry_3(4) := ( pp9(4) and pp10(3) ) or ( pp11(2) and ( pp9(4) xor pp10(3) )) ;
        sigCSA_sum_3(5) := pp9(5) xor pp10(4) xor pp11(3) ;
        sigCSA_cry_3(5) := ( pp9(5) and pp10(4) ) or ( pp11(3) and ( pp9(5) xor pp10(4) )) ;
        sigCSA_sum_3(6) := pp9(6) xor pp10(5) xor pp11(4) ;
        sigCSA_cry_3(6) := ( pp9(6) and pp10(5) ) or ( pp11(4) and ( pp9(6) xor pp10(5) )) ;
        sigCSA_sum_3(7) := pp9(7) xor pp10(6) xor pp11(5) ;
        sigCSA_cry_3(7) := ( pp9(7) and pp10(6) ) or ( pp11(5) and ( pp9(7) xor pp10(6) )) ;
        sigCSA_sum_3(8) := pp9(8) xor pp10(7) xor pp11(6) ;
        sigCSA_cry_3(8) := ( pp9(8) and pp10(7) ) or ( pp11(6) and ( pp9(8) xor pp10(7) )) ;
        sigCSA_sum_3(9) := pp9(9) xor pp10(8) xor pp11(7) ;
        sigCSA_cry_3(9) := ( pp9(9) and pp10(8) ) or ( pp11(7) and ( pp9(9) xor pp10(8) )) ;
        sigCSA_sum_3(10) := pp9(10) xor pp10(9) xor pp11(8) ;
        sigCSA_cry_3(10) := ( pp9(10) and pp10(9) ) or ( pp11(8) and ( pp9(10) xor pp10(9) )) ;
        sigCSA_sum_3(11) := pp9(11) xor pp10(10) xor pp11(9) ;
        sigCSA_cry_3(11) := ( pp9(11) and pp10(10) ) or ( pp11(9) and ( pp9(11) xor pp10(10) )) ;
        sigCSA_sum_3(12) := pp9(12) xor pp10(11) xor pp11(10) ;
        sigCSA_cry_3(12) := ( pp9(12) and pp10(11) ) or ( pp11(10) and ( pp9(12) xor pp10(11) )) ;
        sigCSA_sum_3(13) := pp9(13) xor pp10(12) xor pp11(11) ;
        sigCSA_cry_3(13) := ( pp9(13) and pp10(12) ) or ( pp11(11) and ( pp9(13) xor pp10(12) )) ;
        sigCSA_sum_3(14) := pp9(14) xor pp10(13) xor pp11(12) ;
        sigCSA_cry_3(14) := ( pp9(14) and pp10(13) ) or ( pp11(12) and ( pp9(14) xor pp10(13) )) ;
        sigCSA_sum_3(15) := pp9(15) xor pp10(14) xor pp11(13) ;
        sigCSA_cry_3(15) := ( pp9(15) and pp10(14) ) or ( pp11(13) and ( pp9(15) xor pp10(14) )) ;
        sigCSA_sum_3(16) := '0' xor pp10(15) xor pp11(14) ;
        sigCSA_cry_3(16) := ( '0' and pp10(15) ) or ( pp11(14) and ( '0' xor pp10(15) )) ;
        sigCSA_sum_3(17) := '0' xor '0' xor pp11(15) ;
        sigCSA_cry_3(17) := ( '0' and '0' ) or ( pp11(15) and ( '0' xor '0' )) ;
-- csa : 4
-- generating sigCSA_sum_4 and sigCSA_cry_4

        sigCSA_sum_4(0) := pp12(0) xor '0' xor '0' ;
        sigCSA_cry_4(0) := ( pp12(0) and '0' ) or ( '0' and ( pp12(0) xor '0' )) ;
        sigCSA_sum_4(1) := pp12(1) xor pp13(0) xor '0' ;
        sigCSA_cry_4(1) := ( pp12(1) and pp13(0) ) or ( '0' and ( pp12(1) xor pp13(0) )) ;
        sigCSA_sum_4(2) := pp12(2) xor pp13(1) xor pp14(0) ;
        sigCSA_cry_4(2) := ( pp12(2) and pp13(1) ) or ( pp14(0) and ( pp12(2) xor pp13(1) )) ;
        sigCSA_sum_4(3) := pp12(3) xor pp13(2) xor pp14(1) ;
        sigCSA_cry_4(3) := ( pp12(3) and pp13(2) ) or ( pp14(1) and ( pp12(3) xor pp13(2) )) ;
        sigCSA_sum_4(4) := pp12(4) xor pp13(3) xor pp14(2) ;
        sigCSA_cry_4(4) := ( pp12(4) and pp13(3) ) or ( pp14(2) and ( pp12(4) xor pp13(3) )) ;
        sigCSA_sum_4(5) := pp12(5) xor pp13(4) xor pp14(3) ;
        sigCSA_cry_4(5) := ( pp12(5) and pp13(4) ) or ( pp14(3) and ( pp12(5) xor pp13(4) )) ;
        sigCSA_sum_4(6) := pp12(6) xor pp13(5) xor pp14(4) ;
        sigCSA_cry_4(6) := ( pp12(6) and pp13(5) ) or ( pp14(4) and ( pp12(6) xor pp13(5) )) ;
        sigCSA_sum_4(7) := pp12(7) xor pp13(6) xor pp14(5) ;
        sigCSA_cry_4(7) := ( pp12(7) and pp13(6) ) or ( pp14(5) and ( pp12(7) xor pp13(6) )) ;
        sigCSA_sum_4(8) := pp12(8) xor pp13(7) xor pp14(6) ;
        sigCSA_cry_4(8) := ( pp12(8) and pp13(7) ) or ( pp14(6) and ( pp12(8) xor pp13(7) )) ;
        sigCSA_sum_4(9) := pp12(9) xor pp13(8) xor pp14(7) ;
        sigCSA_cry_4(9) := ( pp12(9) and pp13(8) ) or ( pp14(7) and ( pp12(9) xor pp13(8) )) ;
        sigCSA_sum_4(10) := pp12(10) xor pp13(9) xor pp14(8) ;
        sigCSA_cry_4(10) := ( pp12(10) and pp13(9) ) or ( pp14(8) and ( pp12(10) xor pp13(9) )) ;
        sigCSA_sum_4(11) := pp12(11) xor pp13(10) xor pp14(9) ;
        sigCSA_cry_4(11) := ( pp12(11) and pp13(10) ) or ( pp14(9) and ( pp12(11) xor pp13(10) )) ;
        sigCSA_sum_4(12) := pp12(12) xor pp13(11) xor pp14(10) ;
        sigCSA_cry_4(12) := ( pp12(12) and pp13(11) ) or ( pp14(10) and ( pp12(12) xor pp13(11) )) ;
        sigCSA_sum_4(13) := pp12(13) xor pp13(12) xor pp14(11) ;
        sigCSA_cry_4(13) := ( pp12(13) and pp13(12) ) or ( pp14(11) and ( pp12(13) xor pp13(12) )) ;
        sigCSA_sum_4(14) := pp12(14) xor pp13(13) xor pp14(12) ;
        sigCSA_cry_4(14) := ( pp12(14) and pp13(13) ) or ( pp14(12) and ( pp12(14) xor pp13(13) )) ;
        sigCSA_sum_4(15) := pp12(15) xor pp13(14) xor pp14(13) ;
        sigCSA_cry_4(15) := ( pp12(15) and pp13(14) ) or ( pp14(13) and ( pp12(15) xor pp13(14) )) ;
        sigCSA_sum_4(16) := '0' xor pp13(15) xor pp14(14) ;
        sigCSA_cry_4(16) := ( '0' and pp13(15) ) or ( pp14(14) and ( '0' xor pp13(15) )) ;
        sigCSA_sum_4(17) := '0' xor '0' xor pp14(15) ;
        sigCSA_cry_4(17) := ( '0' and '0' ) or ( pp14(15) and ( '0' xor '0' )) ;
-- csa : 5
-- generating sigCSA_sum_5 and sigCSA_cry_5

        sigCSA_sum_5(0) := sigCSA_sum_0(0) xor '0' xor '0' ;
        sigCSA_cry_5(0) := ( sigCSA_sum_0(0) and '0' ) or ( '0' and ( sigCSA_sum_0(0) xor '0' )) ;
        sigCSA_sum_5(1) := sigCSA_sum_0(1) xor sigCSA_cry_0(0) xor '0' ;
        sigCSA_cry_5(1) := ( sigCSA_sum_0(1) and sigCSA_cry_0(0) ) or ( '0' and ( sigCSA_sum_0(1) xor sigCSA_cry_0(0) )) ;
        sigCSA_sum_5(2) := sigCSA_sum_0(2) xor sigCSA_cry_0(1) xor '0' ;
        sigCSA_cry_5(2) := ( sigCSA_sum_0(2) and sigCSA_cry_0(1) ) or ( '0' and ( sigCSA_sum_0(2) xor sigCSA_cry_0(1) )) ;
        sigCSA_sum_5(3) := sigCSA_sum_0(3) xor sigCSA_cry_0(2) xor sigCSA_sum_1(0) ;
        sigCSA_cry_5(3) := ( sigCSA_sum_0(3) and sigCSA_cry_0(2) ) or ( sigCSA_sum_1(0) and ( sigCSA_sum_0(3) xor sigCSA_cry_0(2) )) ;
        sigCSA_sum_5(4) := sigCSA_sum_0(4) xor sigCSA_cry_0(3) xor sigCSA_sum_1(1) ;
        sigCSA_cry_5(4) := ( sigCSA_sum_0(4) and sigCSA_cry_0(3) ) or ( sigCSA_sum_1(1) and ( sigCSA_sum_0(4) xor sigCSA_cry_0(3) )) ;
        sigCSA_sum_5(5) := sigCSA_sum_0(5) xor sigCSA_cry_0(4) xor sigCSA_sum_1(2) ;
        sigCSA_cry_5(5) := ( sigCSA_sum_0(5) and sigCSA_cry_0(4) ) or ( sigCSA_sum_1(2) and ( sigCSA_sum_0(5) xor sigCSA_cry_0(4) )) ;
        sigCSA_sum_5(6) := sigCSA_sum_0(6) xor sigCSA_cry_0(5) xor sigCSA_sum_1(3) ;
        sigCSA_cry_5(6) := ( sigCSA_sum_0(6) and sigCSA_cry_0(5) ) or ( sigCSA_sum_1(3) and ( sigCSA_sum_0(6) xor sigCSA_cry_0(5) )) ;
        sigCSA_sum_5(7) := sigCSA_sum_0(7) xor sigCSA_cry_0(6) xor sigCSA_sum_1(4) ;
        sigCSA_cry_5(7) := ( sigCSA_sum_0(7) and sigCSA_cry_0(6) ) or ( sigCSA_sum_1(4) and ( sigCSA_sum_0(7) xor sigCSA_cry_0(6) )) ;
        sigCSA_sum_5(8) := sigCSA_sum_0(8) xor sigCSA_cry_0(7) xor sigCSA_sum_1(5) ;
        sigCSA_cry_5(8) := ( sigCSA_sum_0(8) and sigCSA_cry_0(7) ) or ( sigCSA_sum_1(5) and ( sigCSA_sum_0(8) xor sigCSA_cry_0(7) )) ;
        sigCSA_sum_5(9) := sigCSA_sum_0(9) xor sigCSA_cry_0(8) xor sigCSA_sum_1(6) ;
        sigCSA_cry_5(9) := ( sigCSA_sum_0(9) and sigCSA_cry_0(8) ) or ( sigCSA_sum_1(6) and ( sigCSA_sum_0(9) xor sigCSA_cry_0(8) )) ;
        sigCSA_sum_5(10) := sigCSA_sum_0(10) xor sigCSA_cry_0(9) xor sigCSA_sum_1(7) ;
        sigCSA_cry_5(10) := ( sigCSA_sum_0(10) and sigCSA_cry_0(9) ) or ( sigCSA_sum_1(7) and ( sigCSA_sum_0(10) xor sigCSA_cry_0(9) )) ;
        sigCSA_sum_5(11) := sigCSA_sum_0(11) xor sigCSA_cry_0(10) xor sigCSA_sum_1(8) ;
        sigCSA_cry_5(11) := ( sigCSA_sum_0(11) and sigCSA_cry_0(10) ) or ( sigCSA_sum_1(8) and ( sigCSA_sum_0(11) xor sigCSA_cry_0(10) )) ;
        sigCSA_sum_5(12) := sigCSA_sum_0(12) xor sigCSA_cry_0(11) xor sigCSA_sum_1(9) ;
        sigCSA_cry_5(12) := ( sigCSA_sum_0(12) and sigCSA_cry_0(11) ) or ( sigCSA_sum_1(9) and ( sigCSA_sum_0(12) xor sigCSA_cry_0(11) )) ;
        sigCSA_sum_5(13) := sigCSA_sum_0(13) xor sigCSA_cry_0(12) xor sigCSA_sum_1(10) ;
        sigCSA_cry_5(13) := ( sigCSA_sum_0(13) and sigCSA_cry_0(12) ) or ( sigCSA_sum_1(10) and ( sigCSA_sum_0(13) xor sigCSA_cry_0(12) )) ;
        sigCSA_sum_5(14) := sigCSA_sum_0(14) xor sigCSA_cry_0(13) xor sigCSA_sum_1(11) ;
        sigCSA_cry_5(14) := ( sigCSA_sum_0(14) and sigCSA_cry_0(13) ) or ( sigCSA_sum_1(11) and ( sigCSA_sum_0(14) xor sigCSA_cry_0(13) )) ;
        sigCSA_sum_5(15) := sigCSA_sum_0(15) xor sigCSA_cry_0(14) xor sigCSA_sum_1(12) ;
        sigCSA_cry_5(15) := ( sigCSA_sum_0(15) and sigCSA_cry_0(14) ) or ( sigCSA_sum_1(12) and ( sigCSA_sum_0(15) xor sigCSA_cry_0(14) )) ;
        sigCSA_sum_5(16) := sigCSA_sum_0(16) xor sigCSA_cry_0(15) xor sigCSA_sum_1(13) ;
        sigCSA_cry_5(16) := ( sigCSA_sum_0(16) and sigCSA_cry_0(15) ) or ( sigCSA_sum_1(13) and ( sigCSA_sum_0(16) xor sigCSA_cry_0(15) )) ;
        sigCSA_sum_5(17) := sigCSA_sum_0(17) xor sigCSA_cry_0(16) xor sigCSA_sum_1(14) ;
        sigCSA_cry_5(17) := ( sigCSA_sum_0(17) and sigCSA_cry_0(16) ) or ( sigCSA_sum_1(14) and ( sigCSA_sum_0(17) xor sigCSA_cry_0(16) )) ;
        sigCSA_sum_5(18) := '0' xor sigCSA_cry_0(17) xor sigCSA_sum_1(15) ;
        sigCSA_cry_5(18) := ( '0' and sigCSA_cry_0(17) ) or ( sigCSA_sum_1(15) and ( '0' xor sigCSA_cry_0(17) )) ;
        sigCSA_sum_5(19) := '0' xor '0' xor sigCSA_sum_1(16) ;
        sigCSA_cry_5(19) := ( '0' and '0' ) or ( sigCSA_sum_1(16) and ( '0' xor '0' )) ;
        sigCSA_sum_5(20) := '0' xor '0' xor sigCSA_sum_1(17) ;
        sigCSA_cry_5(20) := ( '0' and '0' ) or ( sigCSA_sum_1(17) and ( '0' xor '0' )) ;
-- csa : 6
-- generating sigCSA_sum_6 and sigCSA_cry_6

        sigCSA_sum_6(0) := sigCSA_cry_1(0) xor '0' xor '0' ;
        sigCSA_cry_6(0) := ( sigCSA_cry_1(0) and '0' ) or ( '0' and ( sigCSA_cry_1(0) xor '0' )) ;
        sigCSA_sum_6(1) := sigCSA_cry_1(1) xor '0' xor '0' ;
        sigCSA_cry_6(1) := ( sigCSA_cry_1(1) and '0' ) or ( '0' and ( sigCSA_cry_1(1) xor '0' )) ;
        sigCSA_sum_6(2) := sigCSA_cry_1(2) xor sigCSA_sum_2(0) xor '0' ;
        sigCSA_cry_6(2) := ( sigCSA_cry_1(2) and sigCSA_sum_2(0) ) or ( '0' and ( sigCSA_cry_1(2) xor sigCSA_sum_2(0) )) ;
        sigCSA_sum_6(3) := sigCSA_cry_1(3) xor sigCSA_sum_2(1) xor sigCSA_cry_2(0) ;
        sigCSA_cry_6(3) := ( sigCSA_cry_1(3) and sigCSA_sum_2(1) ) or ( sigCSA_cry_2(0) and ( sigCSA_cry_1(3) xor sigCSA_sum_2(1) )) ;
        sigCSA_sum_6(4) := sigCSA_cry_1(4) xor sigCSA_sum_2(2) xor sigCSA_cry_2(1) ;
        sigCSA_cry_6(4) := ( sigCSA_cry_1(4) and sigCSA_sum_2(2) ) or ( sigCSA_cry_2(1) and ( sigCSA_cry_1(4) xor sigCSA_sum_2(2) )) ;
        sigCSA_sum_6(5) := sigCSA_cry_1(5) xor sigCSA_sum_2(3) xor sigCSA_cry_2(2) ;
        sigCSA_cry_6(5) := ( sigCSA_cry_1(5) and sigCSA_sum_2(3) ) or ( sigCSA_cry_2(2) and ( sigCSA_cry_1(5) xor sigCSA_sum_2(3) )) ;
        sigCSA_sum_6(6) := sigCSA_cry_1(6) xor sigCSA_sum_2(4) xor sigCSA_cry_2(3) ;
        sigCSA_cry_6(6) := ( sigCSA_cry_1(6) and sigCSA_sum_2(4) ) or ( sigCSA_cry_2(3) and ( sigCSA_cry_1(6) xor sigCSA_sum_2(4) )) ;
        sigCSA_sum_6(7) := sigCSA_cry_1(7) xor sigCSA_sum_2(5) xor sigCSA_cry_2(4) ;
        sigCSA_cry_6(7) := ( sigCSA_cry_1(7) and sigCSA_sum_2(5) ) or ( sigCSA_cry_2(4) and ( sigCSA_cry_1(7) xor sigCSA_sum_2(5) )) ;
        sigCSA_sum_6(8) := sigCSA_cry_1(8) xor sigCSA_sum_2(6) xor sigCSA_cry_2(5) ;
        sigCSA_cry_6(8) := ( sigCSA_cry_1(8) and sigCSA_sum_2(6) ) or ( sigCSA_cry_2(5) and ( sigCSA_cry_1(8) xor sigCSA_sum_2(6) )) ;
        sigCSA_sum_6(9) := sigCSA_cry_1(9) xor sigCSA_sum_2(7) xor sigCSA_cry_2(6) ;
        sigCSA_cry_6(9) := ( sigCSA_cry_1(9) and sigCSA_sum_2(7) ) or ( sigCSA_cry_2(6) and ( sigCSA_cry_1(9) xor sigCSA_sum_2(7) )) ;
        sigCSA_sum_6(10) := sigCSA_cry_1(10) xor sigCSA_sum_2(8) xor sigCSA_cry_2(7) ;
        sigCSA_cry_6(10) := ( sigCSA_cry_1(10) and sigCSA_sum_2(8) ) or ( sigCSA_cry_2(7) and ( sigCSA_cry_1(10) xor sigCSA_sum_2(8) )) ;
        sigCSA_sum_6(11) := sigCSA_cry_1(11) xor sigCSA_sum_2(9) xor sigCSA_cry_2(8) ;
        sigCSA_cry_6(11) := ( sigCSA_cry_1(11) and sigCSA_sum_2(9) ) or ( sigCSA_cry_2(8) and ( sigCSA_cry_1(11) xor sigCSA_sum_2(9) )) ;
        sigCSA_sum_6(12) := sigCSA_cry_1(12) xor sigCSA_sum_2(10) xor sigCSA_cry_2(9) ;
        sigCSA_cry_6(12) := ( sigCSA_cry_1(12) and sigCSA_sum_2(10) ) or ( sigCSA_cry_2(9) and ( sigCSA_cry_1(12) xor sigCSA_sum_2(10) )) ;
        sigCSA_sum_6(13) := sigCSA_cry_1(13) xor sigCSA_sum_2(11) xor sigCSA_cry_2(10) ;
        sigCSA_cry_6(13) := ( sigCSA_cry_1(13) and sigCSA_sum_2(11) ) or ( sigCSA_cry_2(10) and ( sigCSA_cry_1(13) xor sigCSA_sum_2(11) )) ;
        sigCSA_sum_6(14) := sigCSA_cry_1(14) xor sigCSA_sum_2(12) xor sigCSA_cry_2(11) ;
        sigCSA_cry_6(14) := ( sigCSA_cry_1(14) and sigCSA_sum_2(12) ) or ( sigCSA_cry_2(11) and ( sigCSA_cry_1(14) xor sigCSA_sum_2(12) )) ;
        sigCSA_sum_6(15) := sigCSA_cry_1(15) xor sigCSA_sum_2(13) xor sigCSA_cry_2(12) ;
        sigCSA_cry_6(15) := ( sigCSA_cry_1(15) and sigCSA_sum_2(13) ) or ( sigCSA_cry_2(12) and ( sigCSA_cry_1(15) xor sigCSA_sum_2(13) )) ;
        sigCSA_sum_6(16) := sigCSA_cry_1(16) xor sigCSA_sum_2(14) xor sigCSA_cry_2(13) ;
        sigCSA_cry_6(16) := ( sigCSA_cry_1(16) and sigCSA_sum_2(14) ) or ( sigCSA_cry_2(13) and ( sigCSA_cry_1(16) xor sigCSA_sum_2(14) )) ;
        sigCSA_sum_6(17) := sigCSA_cry_1(17) xor sigCSA_sum_2(15) xor sigCSA_cry_2(14) ;
        sigCSA_cry_6(17) := ( sigCSA_cry_1(17) and sigCSA_sum_2(15) ) or ( sigCSA_cry_2(14) and ( sigCSA_cry_1(17) xor sigCSA_sum_2(15) )) ;
        sigCSA_sum_6(18) := '0' xor sigCSA_sum_2(16) xor sigCSA_cry_2(15) ;
        sigCSA_cry_6(18) := ( '0' and sigCSA_sum_2(16) ) or ( sigCSA_cry_2(15) and ( '0' xor sigCSA_sum_2(16) )) ;
        sigCSA_sum_6(19) := '0' xor sigCSA_sum_2(17) xor sigCSA_cry_2(16) ;
        sigCSA_cry_6(19) := ( '0' and sigCSA_sum_2(17) ) or ( sigCSA_cry_2(16) and ( '0' xor sigCSA_sum_2(17) )) ;
        sigCSA_sum_6(20) := '0' xor '0' xor sigCSA_cry_2(17) ;
        sigCSA_cry_6(20) := ( '0' and '0' ) or ( sigCSA_cry_2(17) and ( '0' xor '0' )) ;
-- csa : 7
-- generating sigCSA_sum_7 and sigCSA_cry_7

        sigCSA_sum_7(0) := sigCSA_sum_3(0) xor '0' xor '0' ;
        sigCSA_cry_7(0) := ( sigCSA_sum_3(0) and '0' ) or ( '0' and ( sigCSA_sum_3(0) xor '0' )) ;
        sigCSA_sum_7(1) := sigCSA_sum_3(1) xor sigCSA_cry_3(0) xor '0' ;
        sigCSA_cry_7(1) := ( sigCSA_sum_3(1) and sigCSA_cry_3(0) ) or ( '0' and ( sigCSA_sum_3(1) xor sigCSA_cry_3(0) )) ;
        sigCSA_sum_7(2) := sigCSA_sum_3(2) xor sigCSA_cry_3(1) xor '0' ;
        sigCSA_cry_7(2) := ( sigCSA_sum_3(2) and sigCSA_cry_3(1) ) or ( '0' and ( sigCSA_sum_3(2) xor sigCSA_cry_3(1) )) ;
        sigCSA_sum_7(3) := sigCSA_sum_3(3) xor sigCSA_cry_3(2) xor sigCSA_sum_4(0) ;
        sigCSA_cry_7(3) := ( sigCSA_sum_3(3) and sigCSA_cry_3(2) ) or ( sigCSA_sum_4(0) and ( sigCSA_sum_3(3) xor sigCSA_cry_3(2) )) ;
        sigCSA_sum_7(4) := sigCSA_sum_3(4) xor sigCSA_cry_3(3) xor sigCSA_sum_4(1) ;
        sigCSA_cry_7(4) := ( sigCSA_sum_3(4) and sigCSA_cry_3(3) ) or ( sigCSA_sum_4(1) and ( sigCSA_sum_3(4) xor sigCSA_cry_3(3) )) ;
        sigCSA_sum_7(5) := sigCSA_sum_3(5) xor sigCSA_cry_3(4) xor sigCSA_sum_4(2) ;
        sigCSA_cry_7(5) := ( sigCSA_sum_3(5) and sigCSA_cry_3(4) ) or ( sigCSA_sum_4(2) and ( sigCSA_sum_3(5) xor sigCSA_cry_3(4) )) ;
        sigCSA_sum_7(6) := sigCSA_sum_3(6) xor sigCSA_cry_3(5) xor sigCSA_sum_4(3) ;
        sigCSA_cry_7(6) := ( sigCSA_sum_3(6) and sigCSA_cry_3(5) ) or ( sigCSA_sum_4(3) and ( sigCSA_sum_3(6) xor sigCSA_cry_3(5) )) ;
        sigCSA_sum_7(7) := sigCSA_sum_3(7) xor sigCSA_cry_3(6) xor sigCSA_sum_4(4) ;
        sigCSA_cry_7(7) := ( sigCSA_sum_3(7) and sigCSA_cry_3(6) ) or ( sigCSA_sum_4(4) and ( sigCSA_sum_3(7) xor sigCSA_cry_3(6) )) ;
        sigCSA_sum_7(8) := sigCSA_sum_3(8) xor sigCSA_cry_3(7) xor sigCSA_sum_4(5) ;
        sigCSA_cry_7(8) := ( sigCSA_sum_3(8) and sigCSA_cry_3(7) ) or ( sigCSA_sum_4(5) and ( sigCSA_sum_3(8) xor sigCSA_cry_3(7) )) ;
        sigCSA_sum_7(9) := sigCSA_sum_3(9) xor sigCSA_cry_3(8) xor sigCSA_sum_4(6) ;
        sigCSA_cry_7(9) := ( sigCSA_sum_3(9) and sigCSA_cry_3(8) ) or ( sigCSA_sum_4(6) and ( sigCSA_sum_3(9) xor sigCSA_cry_3(8) )) ;
        sigCSA_sum_7(10) := sigCSA_sum_3(10) xor sigCSA_cry_3(9) xor sigCSA_sum_4(7) ;
        sigCSA_cry_7(10) := ( sigCSA_sum_3(10) and sigCSA_cry_3(9) ) or ( sigCSA_sum_4(7) and ( sigCSA_sum_3(10) xor sigCSA_cry_3(9) )) ;
        sigCSA_sum_7(11) := sigCSA_sum_3(11) xor sigCSA_cry_3(10) xor sigCSA_sum_4(8) ;
        sigCSA_cry_7(11) := ( sigCSA_sum_3(11) and sigCSA_cry_3(10) ) or ( sigCSA_sum_4(8) and ( sigCSA_sum_3(11) xor sigCSA_cry_3(10) )) ;
        sigCSA_sum_7(12) := sigCSA_sum_3(12) xor sigCSA_cry_3(11) xor sigCSA_sum_4(9) ;
        sigCSA_cry_7(12) := ( sigCSA_sum_3(12) and sigCSA_cry_3(11) ) or ( sigCSA_sum_4(9) and ( sigCSA_sum_3(12) xor sigCSA_cry_3(11) )) ;
        sigCSA_sum_7(13) := sigCSA_sum_3(13) xor sigCSA_cry_3(12) xor sigCSA_sum_4(10) ;
        sigCSA_cry_7(13) := ( sigCSA_sum_3(13) and sigCSA_cry_3(12) ) or ( sigCSA_sum_4(10) and ( sigCSA_sum_3(13) xor sigCSA_cry_3(12) )) ;
        sigCSA_sum_7(14) := sigCSA_sum_3(14) xor sigCSA_cry_3(13) xor sigCSA_sum_4(11) ;
        sigCSA_cry_7(14) := ( sigCSA_sum_3(14) and sigCSA_cry_3(13) ) or ( sigCSA_sum_4(11) and ( sigCSA_sum_3(14) xor sigCSA_cry_3(13) )) ;
        sigCSA_sum_7(15) := sigCSA_sum_3(15) xor sigCSA_cry_3(14) xor sigCSA_sum_4(12) ;
        sigCSA_cry_7(15) := ( sigCSA_sum_3(15) and sigCSA_cry_3(14) ) or ( sigCSA_sum_4(12) and ( sigCSA_sum_3(15) xor sigCSA_cry_3(14) )) ;
        sigCSA_sum_7(16) := sigCSA_sum_3(16) xor sigCSA_cry_3(15) xor sigCSA_sum_4(13) ;
        sigCSA_cry_7(16) := ( sigCSA_sum_3(16) and sigCSA_cry_3(15) ) or ( sigCSA_sum_4(13) and ( sigCSA_sum_3(16) xor sigCSA_cry_3(15) )) ;
        sigCSA_sum_7(17) := sigCSA_sum_3(17) xor sigCSA_cry_3(16) xor sigCSA_sum_4(14) ;
        sigCSA_cry_7(17) := ( sigCSA_sum_3(17) and sigCSA_cry_3(16) ) or ( sigCSA_sum_4(14) and ( sigCSA_sum_3(17) xor sigCSA_cry_3(16) )) ;
        sigCSA_sum_7(18) := '0' xor sigCSA_cry_3(17) xor sigCSA_sum_4(15) ;
        sigCSA_cry_7(18) := ( '0' and sigCSA_cry_3(17) ) or ( sigCSA_sum_4(15) and ( '0' xor sigCSA_cry_3(17) )) ;
        sigCSA_sum_7(19) := '0' xor '0' xor sigCSA_sum_4(16) ;
        sigCSA_cry_7(19) := ( '0' and '0' ) or ( sigCSA_sum_4(16) and ( '0' xor '0' )) ;
        sigCSA_sum_7(20) := '0' xor '0' xor sigCSA_sum_4(17) ;
        sigCSA_cry_7(20) := ( '0' and '0' ) or ( sigCSA_sum_4(17) and ( '0' xor '0' )) ;
-- csa : 8
-- generating sigCSA_sum_8 and sigCSA_cry_8

        sigCSA_sum_8(0) := sigCSA_sum_5(0) xor '0' xor '0' ;
        sigCSA_cry_8(0) := ( sigCSA_sum_5(0) and '0' ) or ( '0' and ( sigCSA_sum_5(0) xor '0' )) ;
        sigCSA_sum_8(1) := sigCSA_sum_5(1) xor sigCSA_cry_5(0) xor '0' ;
        sigCSA_cry_8(1) := ( sigCSA_sum_5(1) and sigCSA_cry_5(0) ) or ( '0' and ( sigCSA_sum_5(1) xor sigCSA_cry_5(0) )) ;
        sigCSA_sum_8(2) := sigCSA_sum_5(2) xor sigCSA_cry_5(1) xor '0' ;
        sigCSA_cry_8(2) := ( sigCSA_sum_5(2) and sigCSA_cry_5(1) ) or ( '0' and ( sigCSA_sum_5(2) xor sigCSA_cry_5(1) )) ;
        sigCSA_sum_8(3) := sigCSA_sum_5(3) xor sigCSA_cry_5(2) xor '0' ;
        sigCSA_cry_8(3) := ( sigCSA_sum_5(3) and sigCSA_cry_5(2) ) or ( '0' and ( sigCSA_sum_5(3) xor sigCSA_cry_5(2) )) ;
        sigCSA_sum_8(4) := sigCSA_sum_5(4) xor sigCSA_cry_5(3) xor sigCSA_sum_6(0) ;
        sigCSA_cry_8(4) := ( sigCSA_sum_5(4) and sigCSA_cry_5(3) ) or ( sigCSA_sum_6(0) and ( sigCSA_sum_5(4) xor sigCSA_cry_5(3) )) ;
        sigCSA_sum_8(5) := sigCSA_sum_5(5) xor sigCSA_cry_5(4) xor sigCSA_sum_6(1) ;
        sigCSA_cry_8(5) := ( sigCSA_sum_5(5) and sigCSA_cry_5(4) ) or ( sigCSA_sum_6(1) and ( sigCSA_sum_5(5) xor sigCSA_cry_5(4) )) ;
        sigCSA_sum_8(6) := sigCSA_sum_5(6) xor sigCSA_cry_5(5) xor sigCSA_sum_6(2) ;
        sigCSA_cry_8(6) := ( sigCSA_sum_5(6) and sigCSA_cry_5(5) ) or ( sigCSA_sum_6(2) and ( sigCSA_sum_5(6) xor sigCSA_cry_5(5) )) ;
        sigCSA_sum_8(7) := sigCSA_sum_5(7) xor sigCSA_cry_5(6) xor sigCSA_sum_6(3) ;
        sigCSA_cry_8(7) := ( sigCSA_sum_5(7) and sigCSA_cry_5(6) ) or ( sigCSA_sum_6(3) and ( sigCSA_sum_5(7) xor sigCSA_cry_5(6) )) ;
        sigCSA_sum_8(8) := sigCSA_sum_5(8) xor sigCSA_cry_5(7) xor sigCSA_sum_6(4) ;
        sigCSA_cry_8(8) := ( sigCSA_sum_5(8) and sigCSA_cry_5(7) ) or ( sigCSA_sum_6(4) and ( sigCSA_sum_5(8) xor sigCSA_cry_5(7) )) ;
        sigCSA_sum_8(9) := sigCSA_sum_5(9) xor sigCSA_cry_5(8) xor sigCSA_sum_6(5) ;
        sigCSA_cry_8(9) := ( sigCSA_sum_5(9) and sigCSA_cry_5(8) ) or ( sigCSA_sum_6(5) and ( sigCSA_sum_5(9) xor sigCSA_cry_5(8) )) ;
        sigCSA_sum_8(10) := sigCSA_sum_5(10) xor sigCSA_cry_5(9) xor sigCSA_sum_6(6) ;
        sigCSA_cry_8(10) := ( sigCSA_sum_5(10) and sigCSA_cry_5(9) ) or ( sigCSA_sum_6(6) and ( sigCSA_sum_5(10) xor sigCSA_cry_5(9) )) ;
        sigCSA_sum_8(11) := sigCSA_sum_5(11) xor sigCSA_cry_5(10) xor sigCSA_sum_6(7) ;
        sigCSA_cry_8(11) := ( sigCSA_sum_5(11) and sigCSA_cry_5(10) ) or ( sigCSA_sum_6(7) and ( sigCSA_sum_5(11) xor sigCSA_cry_5(10) )) ;
        sigCSA_sum_8(12) := sigCSA_sum_5(12) xor sigCSA_cry_5(11) xor sigCSA_sum_6(8) ;
        sigCSA_cry_8(12) := ( sigCSA_sum_5(12) and sigCSA_cry_5(11) ) or ( sigCSA_sum_6(8) and ( sigCSA_sum_5(12) xor sigCSA_cry_5(11) )) ;
        sigCSA_sum_8(13) := sigCSA_sum_5(13) xor sigCSA_cry_5(12) xor sigCSA_sum_6(9) ;
        sigCSA_cry_8(13) := ( sigCSA_sum_5(13) and sigCSA_cry_5(12) ) or ( sigCSA_sum_6(9) and ( sigCSA_sum_5(13) xor sigCSA_cry_5(12) )) ;
        sigCSA_sum_8(14) := sigCSA_sum_5(14) xor sigCSA_cry_5(13) xor sigCSA_sum_6(10) ;
        sigCSA_cry_8(14) := ( sigCSA_sum_5(14) and sigCSA_cry_5(13) ) or ( sigCSA_sum_6(10) and ( sigCSA_sum_5(14) xor sigCSA_cry_5(13) )) ;
        sigCSA_sum_8(15) := sigCSA_sum_5(15) xor sigCSA_cry_5(14) xor sigCSA_sum_6(11) ;
        sigCSA_cry_8(15) := ( sigCSA_sum_5(15) and sigCSA_cry_5(14) ) or ( sigCSA_sum_6(11) and ( sigCSA_sum_5(15) xor sigCSA_cry_5(14) )) ;
        sigCSA_sum_8(16) := sigCSA_sum_5(16) xor sigCSA_cry_5(15) xor sigCSA_sum_6(12) ;
        sigCSA_cry_8(16) := ( sigCSA_sum_5(16) and sigCSA_cry_5(15) ) or ( sigCSA_sum_6(12) and ( sigCSA_sum_5(16) xor sigCSA_cry_5(15) )) ;
        sigCSA_sum_8(17) := sigCSA_sum_5(17) xor sigCSA_cry_5(16) xor sigCSA_sum_6(13) ;
        sigCSA_cry_8(17) := ( sigCSA_sum_5(17) and sigCSA_cry_5(16) ) or ( sigCSA_sum_6(13) and ( sigCSA_sum_5(17) xor sigCSA_cry_5(16) )) ;
        sigCSA_sum_8(18) := sigCSA_sum_5(18) xor sigCSA_cry_5(17) xor sigCSA_sum_6(14) ;
        sigCSA_cry_8(18) := ( sigCSA_sum_5(18) and sigCSA_cry_5(17) ) or ( sigCSA_sum_6(14) and ( sigCSA_sum_5(18) xor sigCSA_cry_5(17) )) ;
        sigCSA_sum_8(19) := sigCSA_sum_5(19) xor sigCSA_cry_5(18) xor sigCSA_sum_6(15) ;
        sigCSA_cry_8(19) := ( sigCSA_sum_5(19) and sigCSA_cry_5(18) ) or ( sigCSA_sum_6(15) and ( sigCSA_sum_5(19) xor sigCSA_cry_5(18) )) ;
        sigCSA_sum_8(20) := sigCSA_sum_5(20) xor sigCSA_cry_5(19) xor sigCSA_sum_6(16) ;
        sigCSA_cry_8(20) := ( sigCSA_sum_5(20) and sigCSA_cry_5(19) ) or ( sigCSA_sum_6(16) and ( sigCSA_sum_5(20) xor sigCSA_cry_5(19) )) ;
        sigCSA_sum_8(21) := '0' xor sigCSA_cry_5(20) xor sigCSA_sum_6(17) ;
        sigCSA_cry_8(21) := ( '0' and sigCSA_cry_5(20) ) or ( sigCSA_sum_6(17) and ( '0' xor sigCSA_cry_5(20) )) ;
        sigCSA_sum_8(22) := '0' xor '0' xor sigCSA_sum_6(18) ;
        sigCSA_cry_8(22) := ( '0' and '0' ) or ( sigCSA_sum_6(18) and ( '0' xor '0' )) ;
        sigCSA_sum_8(23) := '0' xor '0' xor sigCSA_sum_6(19) ;
        sigCSA_cry_8(23) := ( '0' and '0' ) or ( sigCSA_sum_6(19) and ( '0' xor '0' )) ;
        sigCSA_sum_8(24) := '0' xor '0' xor sigCSA_sum_6(20) ;
        sigCSA_cry_8(24) := ( '0' and '0' ) or ( sigCSA_sum_6(20) and ( '0' xor '0' )) ;
-- csa : 9
-- generating sigCSA_sum_9 and sigCSA_cry_9

        sigCSA_sum_9(0) := sigCSA_cry_6(0) xor '0' xor '0' ;
        sigCSA_cry_9(0) := ( sigCSA_cry_6(0) and '0' ) or ( '0' and ( sigCSA_cry_6(0) xor '0' )) ;
        sigCSA_sum_9(1) := sigCSA_cry_6(1) xor '0' xor '0' ;
        sigCSA_cry_9(1) := ( sigCSA_cry_6(1) and '0' ) or ( '0' and ( sigCSA_cry_6(1) xor '0' )) ;
        sigCSA_sum_9(2) := sigCSA_cry_6(2) xor '0' xor '0' ;
        sigCSA_cry_9(2) := ( sigCSA_cry_6(2) and '0' ) or ( '0' and ( sigCSA_cry_6(2) xor '0' )) ;
        sigCSA_sum_9(3) := sigCSA_cry_6(3) xor '0' xor '0' ;
        sigCSA_cry_9(3) := ( sigCSA_cry_6(3) and '0' ) or ( '0' and ( sigCSA_cry_6(3) xor '0' )) ;
        sigCSA_sum_9(4) := sigCSA_cry_6(4) xor sigCSA_sum_7(0) xor '0' ;
        sigCSA_cry_9(4) := ( sigCSA_cry_6(4) and sigCSA_sum_7(0) ) or ( '0' and ( sigCSA_cry_6(4) xor sigCSA_sum_7(0) )) ;
        sigCSA_sum_9(5) := sigCSA_cry_6(5) xor sigCSA_sum_7(1) xor sigCSA_cry_7(0) ;
        sigCSA_cry_9(5) := ( sigCSA_cry_6(5) and sigCSA_sum_7(1) ) or ( sigCSA_cry_7(0) and ( sigCSA_cry_6(5) xor sigCSA_sum_7(1) )) ;
        sigCSA_sum_9(6) := sigCSA_cry_6(6) xor sigCSA_sum_7(2) xor sigCSA_cry_7(1) ;
        sigCSA_cry_9(6) := ( sigCSA_cry_6(6) and sigCSA_sum_7(2) ) or ( sigCSA_cry_7(1) and ( sigCSA_cry_6(6) xor sigCSA_sum_7(2) )) ;
        sigCSA_sum_9(7) := sigCSA_cry_6(7) xor sigCSA_sum_7(3) xor sigCSA_cry_7(2) ;
        sigCSA_cry_9(7) := ( sigCSA_cry_6(7) and sigCSA_sum_7(3) ) or ( sigCSA_cry_7(2) and ( sigCSA_cry_6(7) xor sigCSA_sum_7(3) )) ;
        sigCSA_sum_9(8) := sigCSA_cry_6(8) xor sigCSA_sum_7(4) xor sigCSA_cry_7(3) ;
        sigCSA_cry_9(8) := ( sigCSA_cry_6(8) and sigCSA_sum_7(4) ) or ( sigCSA_cry_7(3) and ( sigCSA_cry_6(8) xor sigCSA_sum_7(4) )) ;
        sigCSA_sum_9(9) := sigCSA_cry_6(9) xor sigCSA_sum_7(5) xor sigCSA_cry_7(4) ;
        sigCSA_cry_9(9) := ( sigCSA_cry_6(9) and sigCSA_sum_7(5) ) or ( sigCSA_cry_7(4) and ( sigCSA_cry_6(9) xor sigCSA_sum_7(5) )) ;
        sigCSA_sum_9(10) := sigCSA_cry_6(10) xor sigCSA_sum_7(6) xor sigCSA_cry_7(5) ;
        sigCSA_cry_9(10) := ( sigCSA_cry_6(10) and sigCSA_sum_7(6) ) or ( sigCSA_cry_7(5) and ( sigCSA_cry_6(10) xor sigCSA_sum_7(6) )) ;
        sigCSA_sum_9(11) := sigCSA_cry_6(11) xor sigCSA_sum_7(7) xor sigCSA_cry_7(6) ;
        sigCSA_cry_9(11) := ( sigCSA_cry_6(11) and sigCSA_sum_7(7) ) or ( sigCSA_cry_7(6) and ( sigCSA_cry_6(11) xor sigCSA_sum_7(7) )) ;
        sigCSA_sum_9(12) := sigCSA_cry_6(12) xor sigCSA_sum_7(8) xor sigCSA_cry_7(7) ;
        sigCSA_cry_9(12) := ( sigCSA_cry_6(12) and sigCSA_sum_7(8) ) or ( sigCSA_cry_7(7) and ( sigCSA_cry_6(12) xor sigCSA_sum_7(8) )) ;
        sigCSA_sum_9(13) := sigCSA_cry_6(13) xor sigCSA_sum_7(9) xor sigCSA_cry_7(8) ;
        sigCSA_cry_9(13) := ( sigCSA_cry_6(13) and sigCSA_sum_7(9) ) or ( sigCSA_cry_7(8) and ( sigCSA_cry_6(13) xor sigCSA_sum_7(9) )) ;
        sigCSA_sum_9(14) := sigCSA_cry_6(14) xor sigCSA_sum_7(10) xor sigCSA_cry_7(9) ;
        sigCSA_cry_9(14) := ( sigCSA_cry_6(14) and sigCSA_sum_7(10) ) or ( sigCSA_cry_7(9) and ( sigCSA_cry_6(14) xor sigCSA_sum_7(10) )) ;
        sigCSA_sum_9(15) := sigCSA_cry_6(15) xor sigCSA_sum_7(11) xor sigCSA_cry_7(10) ;
        sigCSA_cry_9(15) := ( sigCSA_cry_6(15) and sigCSA_sum_7(11) ) or ( sigCSA_cry_7(10) and ( sigCSA_cry_6(15) xor sigCSA_sum_7(11) )) ;
        sigCSA_sum_9(16) := sigCSA_cry_6(16) xor sigCSA_sum_7(12) xor sigCSA_cry_7(11) ;
        sigCSA_cry_9(16) := ( sigCSA_cry_6(16) and sigCSA_sum_7(12) ) or ( sigCSA_cry_7(11) and ( sigCSA_cry_6(16) xor sigCSA_sum_7(12) )) ;
        sigCSA_sum_9(17) := sigCSA_cry_6(17) xor sigCSA_sum_7(13) xor sigCSA_cry_7(12) ;
        sigCSA_cry_9(17) := ( sigCSA_cry_6(17) and sigCSA_sum_7(13) ) or ( sigCSA_cry_7(12) and ( sigCSA_cry_6(17) xor sigCSA_sum_7(13) )) ;
        sigCSA_sum_9(18) := sigCSA_cry_6(18) xor sigCSA_sum_7(14) xor sigCSA_cry_7(13) ;
        sigCSA_cry_9(18) := ( sigCSA_cry_6(18) and sigCSA_sum_7(14) ) or ( sigCSA_cry_7(13) and ( sigCSA_cry_6(18) xor sigCSA_sum_7(14) )) ;
        sigCSA_sum_9(19) := sigCSA_cry_6(19) xor sigCSA_sum_7(15) xor sigCSA_cry_7(14) ;
        sigCSA_cry_9(19) := ( sigCSA_cry_6(19) and sigCSA_sum_7(15) ) or ( sigCSA_cry_7(14) and ( sigCSA_cry_6(19) xor sigCSA_sum_7(15) )) ;
        sigCSA_sum_9(20) := sigCSA_cry_6(20) xor sigCSA_sum_7(16) xor sigCSA_cry_7(15) ;
        sigCSA_cry_9(20) := ( sigCSA_cry_6(20) and sigCSA_sum_7(16) ) or ( sigCSA_cry_7(15) and ( sigCSA_cry_6(20) xor sigCSA_sum_7(16) )) ;
        sigCSA_sum_9(21) := '0' xor sigCSA_sum_7(17) xor sigCSA_cry_7(16) ;
        sigCSA_cry_9(21) := ( '0' and sigCSA_sum_7(17) ) or ( sigCSA_cry_7(16) and ( '0' xor sigCSA_sum_7(17) )) ;
        sigCSA_sum_9(22) := '0' xor sigCSA_sum_7(18) xor sigCSA_cry_7(17) ;
        sigCSA_cry_9(22) := ( '0' and sigCSA_sum_7(18) ) or ( sigCSA_cry_7(17) and ( '0' xor sigCSA_sum_7(18) )) ;
        sigCSA_sum_9(23) := '0' xor sigCSA_sum_7(19) xor sigCSA_cry_7(18) ;
        sigCSA_cry_9(23) := ( '0' and sigCSA_sum_7(19) ) or ( sigCSA_cry_7(18) and ( '0' xor sigCSA_sum_7(19) )) ;
        sigCSA_sum_9(24) := '0' xor sigCSA_sum_7(20) xor sigCSA_cry_7(19) ;
        sigCSA_cry_9(24) := ( '0' and sigCSA_sum_7(20) ) or ( sigCSA_cry_7(19) and ( '0' xor sigCSA_sum_7(20) )) ;
        sigCSA_sum_9(25) := '0' xor '0' xor sigCSA_cry_7(20) ;
        sigCSA_cry_9(25) := ( '0' and '0' ) or ( sigCSA_cry_7(20) and ( '0' xor '0' )) ;
-- csa : 10
-- generating sigCSA_sum_10 and sigCSA_cry_10

        sigCSA_sum_10(0) := sigCSA_sum_8(0) xor '0' xor '0' ;
        sigCSA_cry_10(0) := ( sigCSA_sum_8(0) and '0' ) or ( '0' and ( sigCSA_sum_8(0) xor '0' )) ;
        sigCSA_sum_10(1) := sigCSA_sum_8(1) xor sigCSA_cry_8(0) xor '0' ;
        sigCSA_cry_10(1) := ( sigCSA_sum_8(1) and sigCSA_cry_8(0) ) or ( '0' and ( sigCSA_sum_8(1) xor sigCSA_cry_8(0) )) ;
        sigCSA_sum_10(2) := sigCSA_sum_8(2) xor sigCSA_cry_8(1) xor '0' ;
        sigCSA_cry_10(2) := ( sigCSA_sum_8(2) and sigCSA_cry_8(1) ) or ( '0' and ( sigCSA_sum_8(2) xor sigCSA_cry_8(1) )) ;
        sigCSA_sum_10(3) := sigCSA_sum_8(3) xor sigCSA_cry_8(2) xor '0' ;
        sigCSA_cry_10(3) := ( sigCSA_sum_8(3) and sigCSA_cry_8(2) ) or ( '0' and ( sigCSA_sum_8(3) xor sigCSA_cry_8(2) )) ;
        sigCSA_sum_10(4) := sigCSA_sum_8(4) xor sigCSA_cry_8(3) xor '0' ;
        sigCSA_cry_10(4) := ( sigCSA_sum_8(4) and sigCSA_cry_8(3) ) or ( '0' and ( sigCSA_sum_8(4) xor sigCSA_cry_8(3) )) ;
        sigCSA_sum_10(5) := sigCSA_sum_8(5) xor sigCSA_cry_8(4) xor sigCSA_sum_9(0) ;
        sigCSA_cry_10(5) := ( sigCSA_sum_8(5) and sigCSA_cry_8(4) ) or ( sigCSA_sum_9(0) and ( sigCSA_sum_8(5) xor sigCSA_cry_8(4) )) ;
        sigCSA_sum_10(6) := sigCSA_sum_8(6) xor sigCSA_cry_8(5) xor sigCSA_sum_9(1) ;
        sigCSA_cry_10(6) := ( sigCSA_sum_8(6) and sigCSA_cry_8(5) ) or ( sigCSA_sum_9(1) and ( sigCSA_sum_8(6) xor sigCSA_cry_8(5) )) ;
        sigCSA_sum_10(7) := sigCSA_sum_8(7) xor sigCSA_cry_8(6) xor sigCSA_sum_9(2) ;
        sigCSA_cry_10(7) := ( sigCSA_sum_8(7) and sigCSA_cry_8(6) ) or ( sigCSA_sum_9(2) and ( sigCSA_sum_8(7) xor sigCSA_cry_8(6) )) ;
        sigCSA_sum_10(8) := sigCSA_sum_8(8) xor sigCSA_cry_8(7) xor sigCSA_sum_9(3) ;
        sigCSA_cry_10(8) := ( sigCSA_sum_8(8) and sigCSA_cry_8(7) ) or ( sigCSA_sum_9(3) and ( sigCSA_sum_8(8) xor sigCSA_cry_8(7) )) ;
        sigCSA_sum_10(9) := sigCSA_sum_8(9) xor sigCSA_cry_8(8) xor sigCSA_sum_9(4) ;
        sigCSA_cry_10(9) := ( sigCSA_sum_8(9) and sigCSA_cry_8(8) ) or ( sigCSA_sum_9(4) and ( sigCSA_sum_8(9) xor sigCSA_cry_8(8) )) ;
        sigCSA_sum_10(10) := sigCSA_sum_8(10) xor sigCSA_cry_8(9) xor sigCSA_sum_9(5) ;
        sigCSA_cry_10(10) := ( sigCSA_sum_8(10) and sigCSA_cry_8(9) ) or ( sigCSA_sum_9(5) and ( sigCSA_sum_8(10) xor sigCSA_cry_8(9) )) ;
        sigCSA_sum_10(11) := sigCSA_sum_8(11) xor sigCSA_cry_8(10) xor sigCSA_sum_9(6) ;
        sigCSA_cry_10(11) := ( sigCSA_sum_8(11) and sigCSA_cry_8(10) ) or ( sigCSA_sum_9(6) and ( sigCSA_sum_8(11) xor sigCSA_cry_8(10) )) ;
        sigCSA_sum_10(12) := sigCSA_sum_8(12) xor sigCSA_cry_8(11) xor sigCSA_sum_9(7) ;
        sigCSA_cry_10(12) := ( sigCSA_sum_8(12) and sigCSA_cry_8(11) ) or ( sigCSA_sum_9(7) and ( sigCSA_sum_8(12) xor sigCSA_cry_8(11) )) ;
        sigCSA_sum_10(13) := sigCSA_sum_8(13) xor sigCSA_cry_8(12) xor sigCSA_sum_9(8) ;
        sigCSA_cry_10(13) := ( sigCSA_sum_8(13) and sigCSA_cry_8(12) ) or ( sigCSA_sum_9(8) and ( sigCSA_sum_8(13) xor sigCSA_cry_8(12) )) ;
        sigCSA_sum_10(14) := sigCSA_sum_8(14) xor sigCSA_cry_8(13) xor sigCSA_sum_9(9) ;
        sigCSA_cry_10(14) := ( sigCSA_sum_8(14) and sigCSA_cry_8(13) ) or ( sigCSA_sum_9(9) and ( sigCSA_sum_8(14) xor sigCSA_cry_8(13) )) ;
        sigCSA_sum_10(15) := sigCSA_sum_8(15) xor sigCSA_cry_8(14) xor sigCSA_sum_9(10) ;
        sigCSA_cry_10(15) := ( sigCSA_sum_8(15) and sigCSA_cry_8(14) ) or ( sigCSA_sum_9(10) and ( sigCSA_sum_8(15) xor sigCSA_cry_8(14) )) ;
        sigCSA_sum_10(16) := sigCSA_sum_8(16) xor sigCSA_cry_8(15) xor sigCSA_sum_9(11) ;
        sigCSA_cry_10(16) := ( sigCSA_sum_8(16) and sigCSA_cry_8(15) ) or ( sigCSA_sum_9(11) and ( sigCSA_sum_8(16) xor sigCSA_cry_8(15) )) ;
        sigCSA_sum_10(17) := sigCSA_sum_8(17) xor sigCSA_cry_8(16) xor sigCSA_sum_9(12) ;
        sigCSA_cry_10(17) := ( sigCSA_sum_8(17) and sigCSA_cry_8(16) ) or ( sigCSA_sum_9(12) and ( sigCSA_sum_8(17) xor sigCSA_cry_8(16) )) ;
        sigCSA_sum_10(18) := sigCSA_sum_8(18) xor sigCSA_cry_8(17) xor sigCSA_sum_9(13) ;
        sigCSA_cry_10(18) := ( sigCSA_sum_8(18) and sigCSA_cry_8(17) ) or ( sigCSA_sum_9(13) and ( sigCSA_sum_8(18) xor sigCSA_cry_8(17) )) ;
        sigCSA_sum_10(19) := sigCSA_sum_8(19) xor sigCSA_cry_8(18) xor sigCSA_sum_9(14) ;
        sigCSA_cry_10(19) := ( sigCSA_sum_8(19) and sigCSA_cry_8(18) ) or ( sigCSA_sum_9(14) and ( sigCSA_sum_8(19) xor sigCSA_cry_8(18) )) ;
        sigCSA_sum_10(20) := sigCSA_sum_8(20) xor sigCSA_cry_8(19) xor sigCSA_sum_9(15) ;
        sigCSA_cry_10(20) := ( sigCSA_sum_8(20) and sigCSA_cry_8(19) ) or ( sigCSA_sum_9(15) and ( sigCSA_sum_8(20) xor sigCSA_cry_8(19) )) ;
        sigCSA_sum_10(21) := sigCSA_sum_8(21) xor sigCSA_cry_8(20) xor sigCSA_sum_9(16) ;
        sigCSA_cry_10(21) := ( sigCSA_sum_8(21) and sigCSA_cry_8(20) ) or ( sigCSA_sum_9(16) and ( sigCSA_sum_8(21) xor sigCSA_cry_8(20) )) ;
        sigCSA_sum_10(22) := sigCSA_sum_8(22) xor sigCSA_cry_8(21) xor sigCSA_sum_9(17) ;
        sigCSA_cry_10(22) := ( sigCSA_sum_8(22) and sigCSA_cry_8(21) ) or ( sigCSA_sum_9(17) and ( sigCSA_sum_8(22) xor sigCSA_cry_8(21) )) ;
        sigCSA_sum_10(23) := sigCSA_sum_8(23) xor sigCSA_cry_8(22) xor sigCSA_sum_9(18) ;
        sigCSA_cry_10(23) := ( sigCSA_sum_8(23) and sigCSA_cry_8(22) ) or ( sigCSA_sum_9(18) and ( sigCSA_sum_8(23) xor sigCSA_cry_8(22) )) ;
        sigCSA_sum_10(24) := sigCSA_sum_8(24) xor sigCSA_cry_8(23) xor sigCSA_sum_9(19) ;
        sigCSA_cry_10(24) := ( sigCSA_sum_8(24) and sigCSA_cry_8(23) ) or ( sigCSA_sum_9(19) and ( sigCSA_sum_8(24) xor sigCSA_cry_8(23) )) ;
        sigCSA_sum_10(25) := '0' xor sigCSA_cry_8(24) xor sigCSA_sum_9(20) ;
        sigCSA_cry_10(25) := ( '0' and sigCSA_cry_8(24) ) or ( sigCSA_sum_9(20) and ( '0' xor sigCSA_cry_8(24) )) ;
        sigCSA_sum_10(26) := '0' xor '0' xor sigCSA_sum_9(21) ;
        sigCSA_cry_10(26) := ( '0' and '0' ) or ( sigCSA_sum_9(21) and ( '0' xor '0' )) ;
        sigCSA_sum_10(27) := '0' xor '0' xor sigCSA_sum_9(22) ;
        sigCSA_cry_10(27) := ( '0' and '0' ) or ( sigCSA_sum_9(22) and ( '0' xor '0' )) ;
        sigCSA_sum_10(28) := '0' xor '0' xor sigCSA_sum_9(23) ;
        sigCSA_cry_10(28) := ( '0' and '0' ) or ( sigCSA_sum_9(23) and ( '0' xor '0' )) ;
        sigCSA_sum_10(29) := '0' xor '0' xor sigCSA_sum_9(24) ;
        sigCSA_cry_10(29) := ( '0' and '0' ) or ( sigCSA_sum_9(24) and ( '0' xor '0' )) ;
        sigCSA_sum_10(30) := '0' xor '0' xor sigCSA_sum_9(25) ;
        sigCSA_cry_10(30) := ( '0' and '0' ) or ( sigCSA_sum_9(25) and ( '0' xor '0' )) ;
-- csa : 11
-- generating sigCSA_sum_11 and sigCSA_cry_11

        sigCSA_sum_11(0) := sigCSA_cry_9(0) xor '0' xor '0' ;
        sigCSA_cry_11(0) := ( sigCSA_cry_9(0) and '0' ) or ( '0' and ( sigCSA_cry_9(0) xor '0' )) ;
        sigCSA_sum_11(1) := sigCSA_cry_9(1) xor '0' xor '0' ;
        sigCSA_cry_11(1) := ( sigCSA_cry_9(1) and '0' ) or ( '0' and ( sigCSA_cry_9(1) xor '0' )) ;
        sigCSA_sum_11(2) := sigCSA_cry_9(2) xor '0' xor '0' ;
        sigCSA_cry_11(2) := ( sigCSA_cry_9(2) and '0' ) or ( '0' and ( sigCSA_cry_9(2) xor '0' )) ;
        sigCSA_sum_11(3) := sigCSA_cry_9(3) xor '0' xor '0' ;
        sigCSA_cry_11(3) := ( sigCSA_cry_9(3) and '0' ) or ( '0' and ( sigCSA_cry_9(3) xor '0' )) ;
        sigCSA_sum_11(4) := sigCSA_cry_9(4) xor '0' xor '0' ;
        sigCSA_cry_11(4) := ( sigCSA_cry_9(4) and '0' ) or ( '0' and ( sigCSA_cry_9(4) xor '0' )) ;
        sigCSA_sum_11(5) := sigCSA_cry_9(5) xor '0' xor '0' ;
        sigCSA_cry_11(5) := ( sigCSA_cry_9(5) and '0' ) or ( '0' and ( sigCSA_cry_9(5) xor '0' )) ;
        sigCSA_sum_11(6) := sigCSA_cry_9(6) xor '0' xor '0' ;
        sigCSA_cry_11(6) := ( sigCSA_cry_9(6) and '0' ) or ( '0' and ( sigCSA_cry_9(6) xor '0' )) ;
        sigCSA_sum_11(7) := sigCSA_cry_9(7) xor sigCSA_cry_4(0) xor '0' ;
        sigCSA_cry_11(7) := ( sigCSA_cry_9(7) and sigCSA_cry_4(0) ) or ( '0' and ( sigCSA_cry_9(7) xor sigCSA_cry_4(0) )) ;
        sigCSA_sum_11(8) := sigCSA_cry_9(8) xor sigCSA_cry_4(1) xor '0' ;
        sigCSA_cry_11(8) := ( sigCSA_cry_9(8) and sigCSA_cry_4(1) ) or ( '0' and ( sigCSA_cry_9(8) xor sigCSA_cry_4(1) )) ;
        sigCSA_sum_11(9) := sigCSA_cry_9(9) xor sigCSA_cry_4(2) xor pp15(0) ;
        sigCSA_cry_11(9) := ( sigCSA_cry_9(9) and sigCSA_cry_4(2) ) or ( pp15(0) and ( sigCSA_cry_9(9) xor sigCSA_cry_4(2) )) ;
        sigCSA_sum_11(10) := sigCSA_cry_9(10) xor sigCSA_cry_4(3) xor pp15(1) ;
        sigCSA_cry_11(10) := ( sigCSA_cry_9(10) and sigCSA_cry_4(3) ) or ( pp15(1) and ( sigCSA_cry_9(10) xor sigCSA_cry_4(3) )) ;
        sigCSA_sum_11(11) := sigCSA_cry_9(11) xor sigCSA_cry_4(4) xor pp15(2) ;
        sigCSA_cry_11(11) := ( sigCSA_cry_9(11) and sigCSA_cry_4(4) ) or ( pp15(2) and ( sigCSA_cry_9(11) xor sigCSA_cry_4(4) )) ;
        sigCSA_sum_11(12) := sigCSA_cry_9(12) xor sigCSA_cry_4(5) xor pp15(3) ;
        sigCSA_cry_11(12) := ( sigCSA_cry_9(12) and sigCSA_cry_4(5) ) or ( pp15(3) and ( sigCSA_cry_9(12) xor sigCSA_cry_4(5) )) ;
        sigCSA_sum_11(13) := sigCSA_cry_9(13) xor sigCSA_cry_4(6) xor pp15(4) ;
        sigCSA_cry_11(13) := ( sigCSA_cry_9(13) and sigCSA_cry_4(6) ) or ( pp15(4) and ( sigCSA_cry_9(13) xor sigCSA_cry_4(6) )) ;
        sigCSA_sum_11(14) := sigCSA_cry_9(14) xor sigCSA_cry_4(7) xor pp15(5) ;
        sigCSA_cry_11(14) := ( sigCSA_cry_9(14) and sigCSA_cry_4(7) ) or ( pp15(5) and ( sigCSA_cry_9(14) xor sigCSA_cry_4(7) )) ;
        sigCSA_sum_11(15) := sigCSA_cry_9(15) xor sigCSA_cry_4(8) xor pp15(6) ;
        sigCSA_cry_11(15) := ( sigCSA_cry_9(15) and sigCSA_cry_4(8) ) or ( pp15(6) and ( sigCSA_cry_9(15) xor sigCSA_cry_4(8) )) ;
        sigCSA_sum_11(16) := sigCSA_cry_9(16) xor sigCSA_cry_4(9) xor pp15(7) ;
        sigCSA_cry_11(16) := ( sigCSA_cry_9(16) and sigCSA_cry_4(9) ) or ( pp15(7) and ( sigCSA_cry_9(16) xor sigCSA_cry_4(9) )) ;
        sigCSA_sum_11(17) := sigCSA_cry_9(17) xor sigCSA_cry_4(10) xor pp15(8) ;
        sigCSA_cry_11(17) := ( sigCSA_cry_9(17) and sigCSA_cry_4(10) ) or ( pp15(8) and ( sigCSA_cry_9(17) xor sigCSA_cry_4(10) )) ;
        sigCSA_sum_11(18) := sigCSA_cry_9(18) xor sigCSA_cry_4(11) xor pp15(9) ;
        sigCSA_cry_11(18) := ( sigCSA_cry_9(18) and sigCSA_cry_4(11) ) or ( pp15(9) and ( sigCSA_cry_9(18) xor sigCSA_cry_4(11) )) ;
        sigCSA_sum_11(19) := sigCSA_cry_9(19) xor sigCSA_cry_4(12) xor pp15(10) ;
        sigCSA_cry_11(19) := ( sigCSA_cry_9(19) and sigCSA_cry_4(12) ) or ( pp15(10) and ( sigCSA_cry_9(19) xor sigCSA_cry_4(12) )) ;
        sigCSA_sum_11(20) := sigCSA_cry_9(20) xor sigCSA_cry_4(13) xor pp15(11) ;
        sigCSA_cry_11(20) := ( sigCSA_cry_9(20) and sigCSA_cry_4(13) ) or ( pp15(11) and ( sigCSA_cry_9(20) xor sigCSA_cry_4(13) )) ;
        sigCSA_sum_11(21) := sigCSA_cry_9(21) xor sigCSA_cry_4(14) xor pp15(12) ;
        sigCSA_cry_11(21) := ( sigCSA_cry_9(21) and sigCSA_cry_4(14) ) or ( pp15(12) and ( sigCSA_cry_9(21) xor sigCSA_cry_4(14) )) ;
        sigCSA_sum_11(22) := sigCSA_cry_9(22) xor sigCSA_cry_4(15) xor pp15(13) ;
        sigCSA_cry_11(22) := ( sigCSA_cry_9(22) and sigCSA_cry_4(15) ) or ( pp15(13) and ( sigCSA_cry_9(22) xor sigCSA_cry_4(15) )) ;
        sigCSA_sum_11(23) := sigCSA_cry_9(23) xor sigCSA_cry_4(16) xor pp15(14) ;
        sigCSA_cry_11(23) := ( sigCSA_cry_9(23) and sigCSA_cry_4(16) ) or ( pp15(14) and ( sigCSA_cry_9(23) xor sigCSA_cry_4(16) )) ;
        sigCSA_sum_11(24) := sigCSA_cry_9(24) xor sigCSA_cry_4(17) xor pp15(15) ;
        sigCSA_cry_11(24) := ( sigCSA_cry_9(24) and sigCSA_cry_4(17) ) or ( pp15(15) and ( sigCSA_cry_9(24) xor sigCSA_cry_4(17) )) ;
        sigCSA_sum_11(25) := sigCSA_cry_9(25) xor '0' xor '0' ;
        sigCSA_cry_11(25) := ( sigCSA_cry_9(25) and '0' ) or ( '0' and ( sigCSA_cry_9(25) xor '0' )) ;
        sigCSA_sum_11(26) := '0' xor '0' xor '0' ;
        sigCSA_cry_11(26) := ( '0' and '0' ) or ( '0' and ( '0' xor '0' )) ;
        sigCSA_sum_11(27) := '0' xor '0' xor '0' ;
        sigCSA_cry_11(27) := ( '0' and '0' ) or ( '0' and ( '0' xor '0' )) ;
        sigCSA_sum_11(28) := '0' xor '0' xor '0' ;
        sigCSA_cry_11(28) := ( '0' and '0' ) or ( '0' and ( '0' xor '0' )) ;
        sigCSA_sum_11(29) := '0' xor '0' xor '0' ;
        sigCSA_cry_11(29) := ( '0' and '0' ) or ( '0' and ( '0' xor '0' )) ;
        sigCSA_sum_11(30) := '0' xor '0' xor '0' ;
        sigCSA_cry_11(30) := ( '0' and '0' ) or ( '0' and ( '0' xor '0' )) ;
-- csa : 12
-- generating sigCSA_sum_12 and sigCSA_cry_12

        sigCSA_sum_12(0) := sigCSA_sum_10(0) xor '0' xor '0' ;
        sigCSA_cry_12(0) := ( sigCSA_sum_10(0) and '0' ) or ( '0' and ( sigCSA_sum_10(0) xor '0' )) ;
        sigCSA_sum_12(1) := sigCSA_sum_10(1) xor sigCSA_cry_10(0) xor '0' ;
        sigCSA_cry_12(1) := ( sigCSA_sum_10(1) and sigCSA_cry_10(0) ) or ( '0' and ( sigCSA_sum_10(1) xor sigCSA_cry_10(0) )) ;
        sigCSA_sum_12(2) := sigCSA_sum_10(2) xor sigCSA_cry_10(1) xor '0' ;
        sigCSA_cry_12(2) := ( sigCSA_sum_10(2) and sigCSA_cry_10(1) ) or ( '0' and ( sigCSA_sum_10(2) xor sigCSA_cry_10(1) )) ;
        sigCSA_sum_12(3) := sigCSA_sum_10(3) xor sigCSA_cry_10(2) xor '0' ;
        sigCSA_cry_12(3) := ( sigCSA_sum_10(3) and sigCSA_cry_10(2) ) or ( '0' and ( sigCSA_sum_10(3) xor sigCSA_cry_10(2) )) ;
        sigCSA_sum_12(4) := sigCSA_sum_10(4) xor sigCSA_cry_10(3) xor '0' ;
        sigCSA_cry_12(4) := ( sigCSA_sum_10(4) and sigCSA_cry_10(3) ) or ( '0' and ( sigCSA_sum_10(4) xor sigCSA_cry_10(3) )) ;
        sigCSA_sum_12(5) := sigCSA_sum_10(5) xor sigCSA_cry_10(4) xor '0' ;
        sigCSA_cry_12(5) := ( sigCSA_sum_10(5) and sigCSA_cry_10(4) ) or ( '0' and ( sigCSA_sum_10(5) xor sigCSA_cry_10(4) )) ;
        sigCSA_sum_12(6) := sigCSA_sum_10(6) xor sigCSA_cry_10(5) xor sigCSA_sum_11(0) ;
        sigCSA_cry_12(6) := ( sigCSA_sum_10(6) and sigCSA_cry_10(5) ) or ( sigCSA_sum_11(0) and ( sigCSA_sum_10(6) xor sigCSA_cry_10(5) )) ;
        sigCSA_sum_12(7) := sigCSA_sum_10(7) xor sigCSA_cry_10(6) xor sigCSA_sum_11(1) ;
        sigCSA_cry_12(7) := ( sigCSA_sum_10(7) and sigCSA_cry_10(6) ) or ( sigCSA_sum_11(1) and ( sigCSA_sum_10(7) xor sigCSA_cry_10(6) )) ;
        sigCSA_sum_12(8) := sigCSA_sum_10(8) xor sigCSA_cry_10(7) xor sigCSA_sum_11(2) ;
        sigCSA_cry_12(8) := ( sigCSA_sum_10(8) and sigCSA_cry_10(7) ) or ( sigCSA_sum_11(2) and ( sigCSA_sum_10(8) xor sigCSA_cry_10(7) )) ;
        sigCSA_sum_12(9) := sigCSA_sum_10(9) xor sigCSA_cry_10(8) xor sigCSA_sum_11(3) ;
        sigCSA_cry_12(9) := ( sigCSA_sum_10(9) and sigCSA_cry_10(8) ) or ( sigCSA_sum_11(3) and ( sigCSA_sum_10(9) xor sigCSA_cry_10(8) )) ;
        sigCSA_sum_12(10) := sigCSA_sum_10(10) xor sigCSA_cry_10(9) xor sigCSA_sum_11(4) ;
        sigCSA_cry_12(10) := ( sigCSA_sum_10(10) and sigCSA_cry_10(9) ) or ( sigCSA_sum_11(4) and ( sigCSA_sum_10(10) xor sigCSA_cry_10(9) )) ;
        sigCSA_sum_12(11) := sigCSA_sum_10(11) xor sigCSA_cry_10(10) xor sigCSA_sum_11(5) ;
        sigCSA_cry_12(11) := ( sigCSA_sum_10(11) and sigCSA_cry_10(10) ) or ( sigCSA_sum_11(5) and ( sigCSA_sum_10(11) xor sigCSA_cry_10(10) )) ;
        sigCSA_sum_12(12) := sigCSA_sum_10(12) xor sigCSA_cry_10(11) xor sigCSA_sum_11(6) ;
        sigCSA_cry_12(12) := ( sigCSA_sum_10(12) and sigCSA_cry_10(11) ) or ( sigCSA_sum_11(6) and ( sigCSA_sum_10(12) xor sigCSA_cry_10(11) )) ;
        sigCSA_sum_12(13) := sigCSA_sum_10(13) xor sigCSA_cry_10(12) xor sigCSA_sum_11(7) ;
        sigCSA_cry_12(13) := ( sigCSA_sum_10(13) and sigCSA_cry_10(12) ) or ( sigCSA_sum_11(7) and ( sigCSA_sum_10(13) xor sigCSA_cry_10(12) )) ;
        sigCSA_sum_12(14) := sigCSA_sum_10(14) xor sigCSA_cry_10(13) xor sigCSA_sum_11(8) ;
        sigCSA_cry_12(14) := ( sigCSA_sum_10(14) and sigCSA_cry_10(13) ) or ( sigCSA_sum_11(8) and ( sigCSA_sum_10(14) xor sigCSA_cry_10(13) )) ;
        sigCSA_sum_12(15) := sigCSA_sum_10(15) xor sigCSA_cry_10(14) xor sigCSA_sum_11(9) ;
        sigCSA_cry_12(15) := ( sigCSA_sum_10(15) and sigCSA_cry_10(14) ) or ( sigCSA_sum_11(9) and ( sigCSA_sum_10(15) xor sigCSA_cry_10(14) )) ;
        sigCSA_sum_12(16) := sigCSA_sum_10(16) xor sigCSA_cry_10(15) xor sigCSA_sum_11(10) ;
        sigCSA_cry_12(16) := ( sigCSA_sum_10(16) and sigCSA_cry_10(15) ) or ( sigCSA_sum_11(10) and ( sigCSA_sum_10(16) xor sigCSA_cry_10(15) )) ;
        sigCSA_sum_12(17) := sigCSA_sum_10(17) xor sigCSA_cry_10(16) xor sigCSA_sum_11(11) ;
        sigCSA_cry_12(17) := ( sigCSA_sum_10(17) and sigCSA_cry_10(16) ) or ( sigCSA_sum_11(11) and ( sigCSA_sum_10(17) xor sigCSA_cry_10(16) )) ;
        sigCSA_sum_12(18) := sigCSA_sum_10(18) xor sigCSA_cry_10(17) xor sigCSA_sum_11(12) ;
        sigCSA_cry_12(18) := ( sigCSA_sum_10(18) and sigCSA_cry_10(17) ) or ( sigCSA_sum_11(12) and ( sigCSA_sum_10(18) xor sigCSA_cry_10(17) )) ;
        sigCSA_sum_12(19) := sigCSA_sum_10(19) xor sigCSA_cry_10(18) xor sigCSA_sum_11(13) ;
        sigCSA_cry_12(19) := ( sigCSA_sum_10(19) and sigCSA_cry_10(18) ) or ( sigCSA_sum_11(13) and ( sigCSA_sum_10(19) xor sigCSA_cry_10(18) )) ;
        sigCSA_sum_12(20) := sigCSA_sum_10(20) xor sigCSA_cry_10(19) xor sigCSA_sum_11(14) ;
        sigCSA_cry_12(20) := ( sigCSA_sum_10(20) and sigCSA_cry_10(19) ) or ( sigCSA_sum_11(14) and ( sigCSA_sum_10(20) xor sigCSA_cry_10(19) )) ;
        sigCSA_sum_12(21) := sigCSA_sum_10(21) xor sigCSA_cry_10(20) xor sigCSA_sum_11(15) ;
        sigCSA_cry_12(21) := ( sigCSA_sum_10(21) and sigCSA_cry_10(20) ) or ( sigCSA_sum_11(15) and ( sigCSA_sum_10(21) xor sigCSA_cry_10(20) )) ;
        sigCSA_sum_12(22) := sigCSA_sum_10(22) xor sigCSA_cry_10(21) xor sigCSA_sum_11(16) ;
        sigCSA_cry_12(22) := ( sigCSA_sum_10(22) and sigCSA_cry_10(21) ) or ( sigCSA_sum_11(16) and ( sigCSA_sum_10(22) xor sigCSA_cry_10(21) )) ;
        sigCSA_sum_12(23) := sigCSA_sum_10(23) xor sigCSA_cry_10(22) xor sigCSA_sum_11(17) ;
        sigCSA_cry_12(23) := ( sigCSA_sum_10(23) and sigCSA_cry_10(22) ) or ( sigCSA_sum_11(17) and ( sigCSA_sum_10(23) xor sigCSA_cry_10(22) )) ;
        sigCSA_sum_12(24) := sigCSA_sum_10(24) xor sigCSA_cry_10(23) xor sigCSA_sum_11(18) ;
        sigCSA_cry_12(24) := ( sigCSA_sum_10(24) and sigCSA_cry_10(23) ) or ( sigCSA_sum_11(18) and ( sigCSA_sum_10(24) xor sigCSA_cry_10(23) )) ;
        sigCSA_sum_12(25) := sigCSA_sum_10(25) xor sigCSA_cry_10(24) xor sigCSA_sum_11(19) ;
        sigCSA_cry_12(25) := ( sigCSA_sum_10(25) and sigCSA_cry_10(24) ) or ( sigCSA_sum_11(19) and ( sigCSA_sum_10(25) xor sigCSA_cry_10(24) )) ;
        sigCSA_sum_12(26) := sigCSA_sum_10(26) xor sigCSA_cry_10(25) xor sigCSA_sum_11(20) ;
        sigCSA_cry_12(26) := ( sigCSA_sum_10(26) and sigCSA_cry_10(25) ) or ( sigCSA_sum_11(20) and ( sigCSA_sum_10(26) xor sigCSA_cry_10(25) )) ;
        sigCSA_sum_12(27) := sigCSA_sum_10(27) xor sigCSA_cry_10(26) xor sigCSA_sum_11(21) ;
        sigCSA_cry_12(27) := ( sigCSA_sum_10(27) and sigCSA_cry_10(26) ) or ( sigCSA_sum_11(21) and ( sigCSA_sum_10(27) xor sigCSA_cry_10(26) )) ;
        sigCSA_sum_12(28) := sigCSA_sum_10(28) xor sigCSA_cry_10(27) xor sigCSA_sum_11(22) ;
        sigCSA_cry_12(28) := ( sigCSA_sum_10(28) and sigCSA_cry_10(27) ) or ( sigCSA_sum_11(22) and ( sigCSA_sum_10(28) xor sigCSA_cry_10(27) )) ;
        sigCSA_sum_12(29) := sigCSA_sum_10(29) xor sigCSA_cry_10(28) xor sigCSA_sum_11(23) ;
        sigCSA_cry_12(29) := ( sigCSA_sum_10(29) and sigCSA_cry_10(28) ) or ( sigCSA_sum_11(23) and ( sigCSA_sum_10(29) xor sigCSA_cry_10(28) )) ;
        sigCSA_sum_12(30) := sigCSA_sum_10(30) xor sigCSA_cry_10(29) xor sigCSA_sum_11(24) ;
        sigCSA_cry_12(30) := ( sigCSA_sum_10(30) and sigCSA_cry_10(29) ) or ( sigCSA_sum_11(24) and ( sigCSA_sum_10(30) xor sigCSA_cry_10(29) )) ;
        sigCSA_sum_12(31) := '0' xor sigCSA_cry_10(30) xor sigCSA_sum_11(25) ;
        sigCSA_cry_12(31) := ( '0' and sigCSA_cry_10(30) ) or ( sigCSA_sum_11(25) and ( '0' xor sigCSA_cry_10(30) )) ;
        sigCSA_sum_12(32) := '0' xor '0' xor sigCSA_sum_11(26) ;
        sigCSA_cry_12(32) := ( '0' and '0' ) or ( sigCSA_sum_11(26) and ( '0' xor '0' )) ;
-- csa : 13
-- generating sigCSA_sum_13 and sigCSA_cry_13

        sigCSA_sum_13(0) := sigCSA_sum_12(0) xor '0' xor '0' ;
        sigCSA_cry_13(0) := ( sigCSA_sum_12(0) and '0' ) or ( '0' and ( sigCSA_sum_12(0) xor '0' )) ;
        sigCSA_sum_13(1) := sigCSA_sum_12(1) xor sigCSA_cry_12(0) xor '0' ;
        sigCSA_cry_13(1) := ( sigCSA_sum_12(1) and sigCSA_cry_12(0) ) or ( '0' and ( sigCSA_sum_12(1) xor sigCSA_cry_12(0) )) ;
        sigCSA_sum_13(2) := sigCSA_sum_12(2) xor sigCSA_cry_12(1) xor '0' ;
        sigCSA_cry_13(2) := ( sigCSA_sum_12(2) and sigCSA_cry_12(1) ) or ( '0' and ( sigCSA_sum_12(2) xor sigCSA_cry_12(1) )) ;
        sigCSA_sum_13(3) := sigCSA_sum_12(3) xor sigCSA_cry_12(2) xor '0' ;
        sigCSA_cry_13(3) := ( sigCSA_sum_12(3) and sigCSA_cry_12(2) ) or ( '0' and ( sigCSA_sum_12(3) xor sigCSA_cry_12(2) )) ;
        sigCSA_sum_13(4) := sigCSA_sum_12(4) xor sigCSA_cry_12(3) xor '0' ;
        sigCSA_cry_13(4) := ( sigCSA_sum_12(4) and sigCSA_cry_12(3) ) or ( '0' and ( sigCSA_sum_12(4) xor sigCSA_cry_12(3) )) ;
        sigCSA_sum_13(5) := sigCSA_sum_12(5) xor sigCSA_cry_12(4) xor '0' ;
        sigCSA_cry_13(5) := ( sigCSA_sum_12(5) and sigCSA_cry_12(4) ) or ( '0' and ( sigCSA_sum_12(5) xor sigCSA_cry_12(4) )) ;
        sigCSA_sum_13(6) := sigCSA_sum_12(6) xor sigCSA_cry_12(5) xor '0' ;
        sigCSA_cry_13(6) := ( sigCSA_sum_12(6) and sigCSA_cry_12(5) ) or ( '0' and ( sigCSA_sum_12(6) xor sigCSA_cry_12(5) )) ;
        sigCSA_sum_13(7) := sigCSA_sum_12(7) xor sigCSA_cry_12(6) xor sigCSA_cry_11(0) ;
        sigCSA_cry_13(7) := ( sigCSA_sum_12(7) and sigCSA_cry_12(6) ) or ( sigCSA_cry_11(0) and ( sigCSA_sum_12(7) xor sigCSA_cry_12(6) )) ;
        sigCSA_sum_13(8) := sigCSA_sum_12(8) xor sigCSA_cry_12(7) xor sigCSA_cry_11(1) ;
        sigCSA_cry_13(8) := ( sigCSA_sum_12(8) and sigCSA_cry_12(7) ) or ( sigCSA_cry_11(1) and ( sigCSA_sum_12(8) xor sigCSA_cry_12(7) )) ;
        sigCSA_sum_13(9) := sigCSA_sum_12(9) xor sigCSA_cry_12(8) xor sigCSA_cry_11(2) ;
        sigCSA_cry_13(9) := ( sigCSA_sum_12(9) and sigCSA_cry_12(8) ) or ( sigCSA_cry_11(2) and ( sigCSA_sum_12(9) xor sigCSA_cry_12(8) )) ;
        sigCSA_sum_13(10) := sigCSA_sum_12(10) xor sigCSA_cry_12(9) xor sigCSA_cry_11(3) ;
        sigCSA_cry_13(10) := ( sigCSA_sum_12(10) and sigCSA_cry_12(9) ) or ( sigCSA_cry_11(3) and ( sigCSA_sum_12(10) xor sigCSA_cry_12(9) )) ;
        sigCSA_sum_13(11) := sigCSA_sum_12(11) xor sigCSA_cry_12(10) xor sigCSA_cry_11(4) ;
        sigCSA_cry_13(11) := ( sigCSA_sum_12(11) and sigCSA_cry_12(10) ) or ( sigCSA_cry_11(4) and ( sigCSA_sum_12(11) xor sigCSA_cry_12(10) )) ;
        sigCSA_sum_13(12) := sigCSA_sum_12(12) xor sigCSA_cry_12(11) xor sigCSA_cry_11(5) ;
        sigCSA_cry_13(12) := ( sigCSA_sum_12(12) and sigCSA_cry_12(11) ) or ( sigCSA_cry_11(5) and ( sigCSA_sum_12(12) xor sigCSA_cry_12(11) )) ;
        sigCSA_sum_13(13) := sigCSA_sum_12(13) xor sigCSA_cry_12(12) xor sigCSA_cry_11(6) ;
        sigCSA_cry_13(13) := ( sigCSA_sum_12(13) and sigCSA_cry_12(12) ) or ( sigCSA_cry_11(6) and ( sigCSA_sum_12(13) xor sigCSA_cry_12(12) )) ;
        sigCSA_sum_13(14) := sigCSA_sum_12(14) xor sigCSA_cry_12(13) xor sigCSA_cry_11(7) ;
        sigCSA_cry_13(14) := ( sigCSA_sum_12(14) and sigCSA_cry_12(13) ) or ( sigCSA_cry_11(7) and ( sigCSA_sum_12(14) xor sigCSA_cry_12(13) )) ;
        sigCSA_sum_13(15) := sigCSA_sum_12(15) xor sigCSA_cry_12(14) xor sigCSA_cry_11(8) ;
        sigCSA_cry_13(15) := ( sigCSA_sum_12(15) and sigCSA_cry_12(14) ) or ( sigCSA_cry_11(8) and ( sigCSA_sum_12(15) xor sigCSA_cry_12(14) )) ;
        sigCSA_sum_13(16) := sigCSA_sum_12(16) xor sigCSA_cry_12(15) xor sigCSA_cry_11(9) ;
        sigCSA_cry_13(16) := ( sigCSA_sum_12(16) and sigCSA_cry_12(15) ) or ( sigCSA_cry_11(9) and ( sigCSA_sum_12(16) xor sigCSA_cry_12(15) )) ;
        sigCSA_sum_13(17) := sigCSA_sum_12(17) xor sigCSA_cry_12(16) xor sigCSA_cry_11(10) ;
        sigCSA_cry_13(17) := ( sigCSA_sum_12(17) and sigCSA_cry_12(16) ) or ( sigCSA_cry_11(10) and ( sigCSA_sum_12(17) xor sigCSA_cry_12(16) )) ;
        sigCSA_sum_13(18) := sigCSA_sum_12(18) xor sigCSA_cry_12(17) xor sigCSA_cry_11(11) ;
        sigCSA_cry_13(18) := ( sigCSA_sum_12(18) and sigCSA_cry_12(17) ) or ( sigCSA_cry_11(11) and ( sigCSA_sum_12(18) xor sigCSA_cry_12(17) )) ;
        sigCSA_sum_13(19) := sigCSA_sum_12(19) xor sigCSA_cry_12(18) xor sigCSA_cry_11(12) ;
        sigCSA_cry_13(19) := ( sigCSA_sum_12(19) and sigCSA_cry_12(18) ) or ( sigCSA_cry_11(12) and ( sigCSA_sum_12(19) xor sigCSA_cry_12(18) )) ;
        sigCSA_sum_13(20) := sigCSA_sum_12(20) xor sigCSA_cry_12(19) xor sigCSA_cry_11(13) ;
        sigCSA_cry_13(20) := ( sigCSA_sum_12(20) and sigCSA_cry_12(19) ) or ( sigCSA_cry_11(13) and ( sigCSA_sum_12(20) xor sigCSA_cry_12(19) )) ;
        sigCSA_sum_13(21) := sigCSA_sum_12(21) xor sigCSA_cry_12(20) xor sigCSA_cry_11(14) ;
        sigCSA_cry_13(21) := ( sigCSA_sum_12(21) and sigCSA_cry_12(20) ) or ( sigCSA_cry_11(14) and ( sigCSA_sum_12(21) xor sigCSA_cry_12(20) )) ;
        sigCSA_sum_13(22) := sigCSA_sum_12(22) xor sigCSA_cry_12(21) xor sigCSA_cry_11(15) ;
        sigCSA_cry_13(22) := ( sigCSA_sum_12(22) and sigCSA_cry_12(21) ) or ( sigCSA_cry_11(15) and ( sigCSA_sum_12(22) xor sigCSA_cry_12(21) )) ;
        sigCSA_sum_13(23) := sigCSA_sum_12(23) xor sigCSA_cry_12(22) xor sigCSA_cry_11(16) ;
        sigCSA_cry_13(23) := ( sigCSA_sum_12(23) and sigCSA_cry_12(22) ) or ( sigCSA_cry_11(16) and ( sigCSA_sum_12(23) xor sigCSA_cry_12(22) )) ;
        sigCSA_sum_13(24) := sigCSA_sum_12(24) xor sigCSA_cry_12(23) xor sigCSA_cry_11(17) ;
        sigCSA_cry_13(24) := ( sigCSA_sum_12(24) and sigCSA_cry_12(23) ) or ( sigCSA_cry_11(17) and ( sigCSA_sum_12(24) xor sigCSA_cry_12(23) )) ;
        sigCSA_sum_13(25) := sigCSA_sum_12(25) xor sigCSA_cry_12(24) xor sigCSA_cry_11(18) ;
        sigCSA_cry_13(25) := ( sigCSA_sum_12(25) and sigCSA_cry_12(24) ) or ( sigCSA_cry_11(18) and ( sigCSA_sum_12(25) xor sigCSA_cry_12(24) )) ;
        sigCSA_sum_13(26) := sigCSA_sum_12(26) xor sigCSA_cry_12(25) xor sigCSA_cry_11(19) ;
        sigCSA_cry_13(26) := ( sigCSA_sum_12(26) and sigCSA_cry_12(25) ) or ( sigCSA_cry_11(19) and ( sigCSA_sum_12(26) xor sigCSA_cry_12(25) )) ;
        sigCSA_sum_13(27) := sigCSA_sum_12(27) xor sigCSA_cry_12(26) xor sigCSA_cry_11(20) ;
        sigCSA_cry_13(27) := ( sigCSA_sum_12(27) and sigCSA_cry_12(26) ) or ( sigCSA_cry_11(20) and ( sigCSA_sum_12(27) xor sigCSA_cry_12(26) )) ;
        sigCSA_sum_13(28) := sigCSA_sum_12(28) xor sigCSA_cry_12(27) xor sigCSA_cry_11(21) ;
        sigCSA_cry_13(28) := ( sigCSA_sum_12(28) and sigCSA_cry_12(27) ) or ( sigCSA_cry_11(21) and ( sigCSA_sum_12(28) xor sigCSA_cry_12(27) )) ;
        sigCSA_sum_13(29) := sigCSA_sum_12(29) xor sigCSA_cry_12(28) xor sigCSA_cry_11(22) ;
        sigCSA_cry_13(29) := ( sigCSA_sum_12(29) and sigCSA_cry_12(28) ) or ( sigCSA_cry_11(22) and ( sigCSA_sum_12(29) xor sigCSA_cry_12(28) )) ;
        sigCSA_sum_13(30) := sigCSA_sum_12(30) xor sigCSA_cry_12(29) xor sigCSA_cry_11(23) ;
        sigCSA_cry_13(30) := ( sigCSA_sum_12(30) and sigCSA_cry_12(29) ) or ( sigCSA_cry_11(23) and ( sigCSA_sum_12(30) xor sigCSA_cry_12(29) )) ;
        sigCSA_sum_13(31) := sigCSA_sum_12(31) xor sigCSA_cry_12(30) xor sigCSA_cry_11(24) ;
        sigCSA_cry_13(31) := ( sigCSA_sum_12(31) and sigCSA_cry_12(30) ) or ( sigCSA_cry_11(24) and ( sigCSA_sum_12(31) xor sigCSA_cry_12(30) )) ;
        sigCSA_sum_13(32) := sigCSA_sum_12(32) xor sigCSA_cry_12(31) xor '0' ;
        sigCSA_cry_13(32) := ( sigCSA_sum_12(32) and sigCSA_cry_12(31) ) or ( '0' and ( sigCSA_sum_12(32) xor sigCSA_cry_12(31) )) ;
-- ******************
-- the final output
        result_int(0) := sigCSA_sum_13(0);
        result_int(1) := sigCSA_sum_13(1) xor sigCSA_cry_13(0) xor '0' ;
        carry_rca(0) := sigCSA_sum_13(1) and sigCSA_cry_13(0);
        result_int(2) := sigCSA_sum_13(2) xor sigCSA_cry_13(1) xor carry_rca(0);
        carry_rca(1) := ( sigCSA_sum_13(2) and sigCSA_cry_13(1)) or ( carry_rca(0) and ( sigCSA_sum_13(2) xor sigCSA_cry_13(1)));
        result_int(3) := sigCSA_sum_13(3) xor sigCSA_cry_13(2) xor carry_rca(1);
        carry_rca(2) := ( sigCSA_sum_13(3) and sigCSA_cry_13(2)) or ( carry_rca(1) and ( sigCSA_sum_13(3) xor sigCSA_cry_13(2)));
        result_int(4) := sigCSA_sum_13(4) xor sigCSA_cry_13(3) xor carry_rca(2);
        carry_rca(3) := ( sigCSA_sum_13(4) and sigCSA_cry_13(3)) or ( carry_rca(2) and ( sigCSA_sum_13(4) xor sigCSA_cry_13(3)));
        result_int(5) := sigCSA_sum_13(5) xor sigCSA_cry_13(4) xor carry_rca(3);
        carry_rca(4) := ( sigCSA_sum_13(5) and sigCSA_cry_13(4)) or ( carry_rca(3) and ( sigCSA_sum_13(5) xor sigCSA_cry_13(4)));
        result_int(6) := sigCSA_sum_13(6) xor sigCSA_cry_13(5) xor carry_rca(4);
        carry_rca(5) := ( sigCSA_sum_13(6) and sigCSA_cry_13(5)) or ( carry_rca(4) and ( sigCSA_sum_13(6) xor sigCSA_cry_13(5)));
        result_int(7) := sigCSA_sum_13(7) xor sigCSA_cry_13(6) xor carry_rca(5);
        carry_rca(6) := ( sigCSA_sum_13(7) and sigCSA_cry_13(6)) or ( carry_rca(5) and ( sigCSA_sum_13(7) xor sigCSA_cry_13(6)));
        result_int(8) := sigCSA_sum_13(8) xor sigCSA_cry_13(7) xor carry_rca(6);
        carry_rca(7) := ( sigCSA_sum_13(8) and sigCSA_cry_13(7)) or ( carry_rca(6) and ( sigCSA_sum_13(8) xor sigCSA_cry_13(7)));
        result_int(9) := sigCSA_sum_13(9) xor sigCSA_cry_13(8) xor carry_rca(7);
        carry_rca(8) := ( sigCSA_sum_13(9) and sigCSA_cry_13(8)) or ( carry_rca(7) and ( sigCSA_sum_13(9) xor sigCSA_cry_13(8)));
        result_int(10) := sigCSA_sum_13(10) xor sigCSA_cry_13(9) xor carry_rca(8);
        carry_rca(9) := ( sigCSA_sum_13(10) and sigCSA_cry_13(9)) or ( carry_rca(8) and ( sigCSA_sum_13(10) xor sigCSA_cry_13(9)));
        result_int(11) := sigCSA_sum_13(11) xor sigCSA_cry_13(10) xor carry_rca(9);
        carry_rca(10) := ( sigCSA_sum_13(11) and sigCSA_cry_13(10)) or ( carry_rca(9) and ( sigCSA_sum_13(11) xor sigCSA_cry_13(10)));
        result_int(12) := sigCSA_sum_13(12) xor sigCSA_cry_13(11) xor carry_rca(10);
        carry_rca(11) := ( sigCSA_sum_13(12) and sigCSA_cry_13(11)) or ( carry_rca(10) and ( sigCSA_sum_13(12) xor sigCSA_cry_13(11)));
        result_int(13) := sigCSA_sum_13(13) xor sigCSA_cry_13(12) xor carry_rca(11);
        carry_rca(12) := ( sigCSA_sum_13(13) and sigCSA_cry_13(12)) or ( carry_rca(11) and ( sigCSA_sum_13(13) xor sigCSA_cry_13(12)));
        result_int(14) := sigCSA_sum_13(14) xor sigCSA_cry_13(13) xor carry_rca(12);
        carry_rca(13) := ( sigCSA_sum_13(14) and sigCSA_cry_13(13)) or ( carry_rca(12) and ( sigCSA_sum_13(14) xor sigCSA_cry_13(13)));
        result_int(15) := sigCSA_sum_13(15) xor sigCSA_cry_13(14) xor carry_rca(13);
        carry_rca(14) := ( sigCSA_sum_13(15) and sigCSA_cry_13(14)) or ( carry_rca(13) and ( sigCSA_sum_13(15) xor sigCSA_cry_13(14)));
        result_int(16) := sigCSA_sum_13(16) xor sigCSA_cry_13(15) xor carry_rca(14);
        carry_rca(15) := ( sigCSA_sum_13(16) and sigCSA_cry_13(15)) or ( carry_rca(14) and ( sigCSA_sum_13(16) xor sigCSA_cry_13(15)));
        result_int(17) := sigCSA_sum_13(17) xor sigCSA_cry_13(16) xor carry_rca(15);
        carry_rca(16) := ( sigCSA_sum_13(17) and sigCSA_cry_13(16)) or ( carry_rca(15) and ( sigCSA_sum_13(17) xor sigCSA_cry_13(16)));
        result_int(18) := sigCSA_sum_13(18) xor sigCSA_cry_13(17) xor carry_rca(16);
        carry_rca(17) := ( sigCSA_sum_13(18) and sigCSA_cry_13(17)) or ( carry_rca(16) and ( sigCSA_sum_13(18) xor sigCSA_cry_13(17)));
        result_int(19) := sigCSA_sum_13(19) xor sigCSA_cry_13(18) xor carry_rca(17);
        carry_rca(18) := ( sigCSA_sum_13(19) and sigCSA_cry_13(18)) or ( carry_rca(17) and ( sigCSA_sum_13(19) xor sigCSA_cry_13(18)));
        result_int(20) := sigCSA_sum_13(20) xor sigCSA_cry_13(19) xor carry_rca(18);
        carry_rca(19) := ( sigCSA_sum_13(20) and sigCSA_cry_13(19)) or ( carry_rca(18) and ( sigCSA_sum_13(20) xor sigCSA_cry_13(19)));
        result_int(21) := sigCSA_sum_13(21) xor sigCSA_cry_13(20) xor carry_rca(19);
        carry_rca(20) := ( sigCSA_sum_13(21) and sigCSA_cry_13(20)) or ( carry_rca(19) and ( sigCSA_sum_13(21) xor sigCSA_cry_13(20)));
        result_int(22) := sigCSA_sum_13(22) xor sigCSA_cry_13(21) xor carry_rca(20);
        carry_rca(21) := ( sigCSA_sum_13(22) and sigCSA_cry_13(21)) or ( carry_rca(20) and ( sigCSA_sum_13(22) xor sigCSA_cry_13(21)));
        result_int(23) := sigCSA_sum_13(23) xor sigCSA_cry_13(22) xor carry_rca(21);
        carry_rca(22) := ( sigCSA_sum_13(23) and sigCSA_cry_13(22)) or ( carry_rca(21) and ( sigCSA_sum_13(23) xor sigCSA_cry_13(22)));
        result_int(24) := sigCSA_sum_13(24) xor sigCSA_cry_13(23) xor carry_rca(22);
        carry_rca(23) := ( sigCSA_sum_13(24) and sigCSA_cry_13(23)) or ( carry_rca(22) and ( sigCSA_sum_13(24) xor sigCSA_cry_13(23)));
        result_int(25) := sigCSA_sum_13(25) xor sigCSA_cry_13(24) xor carry_rca(23);
        carry_rca(24) := ( sigCSA_sum_13(25) and sigCSA_cry_13(24)) or ( carry_rca(23) and ( sigCSA_sum_13(25) xor sigCSA_cry_13(24)));
        result_int(26) := sigCSA_sum_13(26) xor sigCSA_cry_13(25) xor carry_rca(24);
        carry_rca(25) := ( sigCSA_sum_13(26) and sigCSA_cry_13(25)) or ( carry_rca(24) and ( sigCSA_sum_13(26) xor sigCSA_cry_13(25)));
        result_int(27) := sigCSA_sum_13(27) xor sigCSA_cry_13(26) xor carry_rca(25);
        carry_rca(26) := ( sigCSA_sum_13(27) and sigCSA_cry_13(26)) or ( carry_rca(25) and ( sigCSA_sum_13(27) xor sigCSA_cry_13(26)));
        result_int(28) := sigCSA_sum_13(28) xor sigCSA_cry_13(27) xor carry_rca(26);
        carry_rca(27) := ( sigCSA_sum_13(28) and sigCSA_cry_13(27)) or ( carry_rca(26) and ( sigCSA_sum_13(28) xor sigCSA_cry_13(27)));
        result_int(29) := sigCSA_sum_13(29) xor sigCSA_cry_13(28) xor carry_rca(27);
        carry_rca(28) := ( sigCSA_sum_13(29) and sigCSA_cry_13(28)) or ( carry_rca(27) and ( sigCSA_sum_13(29) xor sigCSA_cry_13(28)));
        result_int(30) := sigCSA_sum_13(30) xor sigCSA_cry_13(29) xor carry_rca(28);
        carry_rca(29) := ( sigCSA_sum_13(30) and sigCSA_cry_13(29)) or ( carry_rca(28) and ( sigCSA_sum_13(30) xor sigCSA_cry_13(29)));
        result_int(31) := sigCSA_sum_13(31) xor sigCSA_cry_13(30) xor carry_rca(29);
        carry_rca(30) := ( sigCSA_sum_13(31) and sigCSA_cry_13(30)) or ( carry_rca(29) and ( sigCSA_sum_13(31) xor sigCSA_cry_13(30)));
        result_int(32) := sigCSA_sum_13(32) xor sigCSA_cry_13(31) xor carry_rca(30);
        carry_rca(31) := ( sigCSA_sum_13(32) and sigCSA_cry_13(31)) or ( carry_rca(30) and ( sigCSA_sum_13(32) xor sigCSA_cry_13(31)));
        result_int(32) := sigCSA_cry_13(31) xor carry_rca(30);
      
        return result_int;        
        end function mul_func;
        
end package body;
